--Engineer     : Navdeep Dahiya
--Date         : 11/15/2018
--Name of file : block_rom.vhd
--Description  : module ROM as block rom

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity blk_rom_4 is
  port (
	-- input side
	clk	: in std_logic;
	rst	: in std_logic;
	addr	: in integer range 0 to 14999; -- address bits
	--output side
	data_o_1	: out std_logic_vector(7 downto 0);
	data_o_2    : out std_logic_vector(7 downto 0);
	data_o_3    : out std_logic_vector(7 downto 0);
	data_o_4    : out std_logic_vector(7 downto 0)
	);
end blk_rom_4;

architecture arch of blk_rom_4 is

signal addr_1 : integer range 0 to 14999;
signal addr_2 : integer range 0 to 14999;
signal addr_3 : integer range 0 to 14999;
signal addr_4 : integer range 0 to 14999;

type rom_t is array(0 to 14999) of std_logic_vector(7 downto 0);

signal rom : rom_t := (
		"01010001",
		"01100111",
		"01100010",
		"01100110",
		"01100101",
		"01100111",
		"01100110",
		"01100110",
		"01100101",
		"01100100",
		"01100101",
		"01101000",
		"01100101",
		"01100101",
		"01100101",
		"01100110",
		"01100110",
		"01100100",
		"01100011",
		"01100001",
		"01100001",
		"01100001",
		"01011111",
		"01011100",
		"01101110",
		"10010011",
		"10101000",
		"10101010",
		"10001010",
		"01011001",
		"01000101",
		"01000011",
		"01000010",
		"01100001",
		"10000010",
		"01111111",
		"10010001",
		"10100101",
		"10101010",
		"10101011",
		"10101101",
		"10101111",
		"10101111",
		"10101111",
		"10101111",
		"10101111",
		"10101111",
		"10101111",
		"10101110",
		"10101011",
		"10101001",
		"10100101",
		"10100001",
		"10011010",
		"10000101",
		"10001001",
		"10011110",
		"10101010",
		"10100111",
		"10011010",
		"10001001",
		"10000011",
		"10000100",
		"10001001",
		"10001100",
		"10010000",
		"10010010",
		"10010011",
		"10010001",
		"10001110",
		"10001010",
		"10000011",
		"01111100",
		"01110101",
		"01101100",
		"01110110",
		"10001111",
		"10100010",
		"10100110",
		"10101000",
		"10100011",
		"10100010",
		"10100011",
		"10100011",
		"10100011",
		"10100100",
		"10100100",
		"10100101",
		"10100110",
		"10100111",
		"10101001",
		"10101101",
		"10110101",
		"10001111",
		"01000000",
		"01010110",
		"10001100",
		"10011001",
		"10100001",
		"10100111",
		"10100011",
		"01110001",
		"01010010",
		"01010110",
		"01011000",
		"01011011",
		"01011110",
		"01011010",
		"01010001",
		"01101100",
		"01101010",
		"01011101",
		"01011001",
		"01010100",
		"01011000",
		"01100000",
		"01100110",
		"01110111",
		"10000100",
		"10001011",
		"10010001",
		"10010011",
		"10010110",
		"10011011",
		"10100001",
		"10011010",
		"10011001",
		"10011010",
		"10011001",
		"10010010",
		"01110011",
		"01011010",
		"01011111",
		"01100110",
		"01100000",
		"01010001",
		"01100001",
		"01110010",
		"01111000",
		"01111100",
		"01111100",
		"01111111",
		"10000111",
		"10010001",
		"10011100",
		"10011111",
		"10011110",
		"10011101",
		"10011010",
		"10010001",
		"01010110",
		"01110010",
		"01101101",
		"01101111",
		"01101110",
		"01101011",
		"01101001",
		"01101010",
		"01100111",
		"01100111",
		"01101000",
		"01101010",
		"01101100",
		"01101010",
		"01101101",
		"01101101",
		"01101101",
		"01101011",
		"01101010",
		"01101010",
		"01101010",
		"01101001",
		"01100101",
		"01100010",
		"01100011",
		"01110011",
		"10010100",
		"10111001",
		"11001010",
		"10111000",
		"10010100",
		"01110110",
		"01100101",
		"01111100",
		"10010000",
		"10000110",
		"10011010",
		"10111101",
		"11000111",
		"11001010",
		"11001101",
		"11010001",
		"11010100",
		"11010100",
		"11010010",
		"11010000",
		"11001111",
		"11001110",
		"11001101",
		"11001000",
		"10111111",
		"10101101",
		"10011100",
		"10011011",
		"10100101",
		"10110001",
		"11000100",
		"10100101",
		"01110001",
		"01011001",
		"01010011",
		"01010110",
		"01011000",
		"01011010",
		"01011011",
		"01011101",
		"01011110",
		"01100010",
		"01100101",
		"01100100",
		"01100100",
		"01101000",
		"01101010",
		"01101000",
		"10000111",
		"10110110",
		"11000011",
		"11000100",
		"11000110",
		"11001101",
		"11010000",
		"11001110",
		"11001101",
		"11001110",
		"11001111",
		"11001111",
		"11010000",
		"11010000",
		"11001110",
		"11001111",
		"11010001",
		"11010110",
		"11010110",
		"01110110",
		"01000011",
		"01011100",
		"10110001",
		"11000110",
		"10111010",
		"10110011",
		"10100100",
		"10010000",
		"10011000",
		"10010001",
		"10001010",
		"10000101",
		"01101011",
		"01011001",
		"01010011",
		"01010111",
		"01011010",
		"01011101",
		"01011111",
		"01101110",
		"01111100",
		"10000101",
		"10010010",
		"10100010",
		"10101011",
		"10110000",
		"10110111",
		"10111010",
		"10111011",
		"10111011",
		"10111101",
		"11000000",
		"11000001",
		"11000001",
		"11000010",
		"11000000",
		"10110101",
		"10010010",
		"01110101",
		"01110111",
		"01101010",
		"01100011",
		"01110101",
		"10000100",
		"10001011",
		"10001111",
		"10010000",
		"10010100",
		"10011101",
		"10100100",
		"10101110",
		"10110100",
		"10110110",
		"10110011",
		"10110011",
		"10101010",
		"01001110",
		"01101010",
		"01100110",
		"01101001",
		"01101000",
		"01100111",
		"01101001",
		"01101100",
		"01101101",
		"01101110",
		"01101010",
		"01100111",
		"01100110",
		"01100101",
		"01101010",
		"01101010",
		"01101011",
		"01101010",
		"01101101",
		"01101010",
		"01101010",
		"01101100",
		"01101010",
		"01101011",
		"01101000",
		"01100110",
		"01100101",
		"01110100",
		"10011010",
		"10111010",
		"11001001",
		"11001001",
		"11000011",
		"10101111",
		"10001110",
		"10000011",
		"10011000",
		"10110110",
		"11000010",
		"11000111",
		"11001100",
		"11010011",
		"11010110",
		"11011001",
		"11011100",
		"11011011",
		"11011001",
		"11010110",
		"11001101",
		"10111010",
		"10100010",
		"10010101",
		"10100010",
		"10110101",
		"10111110",
		"10110010",
		"10001011",
		"01011011",
		"01010011",
		"01010101",
		"01011001",
		"01011001",
		"01011011",
		"01011100",
		"01011101",
		"01011111",
		"01011110",
		"01011101",
		"01011111",
		"01011101",
		"01011101",
		"01011111",
		"01100000",
		"01100001",
		"01101100",
		"10001010",
		"10101011",
		"11000111",
		"11010000",
		"11010000",
		"11001110",
		"11001101",
		"11001110",
		"11010000",
		"11010000",
		"11010001",
		"11010010",
		"11001111",
		"11001100",
		"11001010",
		"11001010",
		"11001111",
		"10100010",
		"01011111",
		"01110000",
		"10001111",
		"11000010",
		"11001010",
		"11000110",
		"11000010",
		"11000000",
		"10100110",
		"10100111",
		"10110001",
		"10100100",
		"10011110",
		"10101000",
		"10010110",
		"01111000",
		"01010011",
		"01000001",
		"01001101",
		"01100010",
		"10000010",
		"10001110",
		"10011000",
		"10011110",
		"10100110",
		"10101011",
		"10101110",
		"10110010",
		"10110100",
		"10110110",
		"10111000",
		"10111001",
		"10111011",
		"10111101",
		"10111111",
		"11000000",
		"11000000",
		"10111111",
		"10110111",
		"10010011",
		"01110001",
		"01011010",
		"01011011",
		"01110010",
		"01111100",
		"01111010",
		"10000001",
		"10001101",
		"10011010",
		"10100010",
		"10101001",
		"10110000",
		"10110011",
		"10110010",
		"10101101",
		"10101001",
		"10100100",
		"01011000",
		"10000111",
		"10000100",
		"10001000",
		"10001101",
		"10010000",
		"10011000",
		"10100000",
		"10100110",
		"10100111",
		"10100100",
		"10010101",
		"01111000",
		"01011111",
		"01011110",
		"01100100",
		"01100110",
		"01100010",
		"01100010",
		"01100010",
		"01100101",
		"01101000",
		"01101000",
		"01100110",
		"01100111",
		"01100110",
		"01100101",
		"01100011",
		"01100000",
		"01101001",
		"10000011",
		"10011110",
		"10101111",
		"10100010",
		"10000010",
		"01111011",
		"10011100",
		"10111010",
		"11000111",
		"11001000",
		"10111000",
		"10100011",
		"10010000",
		"10001001",
		"10000011",
		"01111111",
		"10000011",
		"10010011",
		"10010111",
		"10010100",
		"10100010",
		"10110110",
		"10110101",
		"10010110",
		"01101011",
		"01011001",
		"01011100",
		"01011100",
		"01011010",
		"01011001",
		"01011011",
		"01011100",
		"01011011",
		"01011101",
		"01011110",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01011111",
		"01100001",
		"01100010",
		"01100010",
		"01100001",
		"01100000",
		"01011110",
		"01011111",
		"01110100",
		"10100001",
		"11001010",
		"11011010",
		"11011001",
		"11010100",
		"11010001",
		"11001111",
		"11010000",
		"11001111",
		"11001011",
		"11000101",
		"10111111",
		"10111010",
		"10010110",
		"01101111",
		"01111010",
		"01111111",
		"10011110",
		"10111111",
		"11010000",
		"11001000",
		"11010011",
		"11000010",
		"10100000",
		"10100011",
		"10101111",
		"10110111",
		"10100111",
		"10101001",
		"10110101",
		"10110101",
		"10100001",
		"01011000",
		"01001101",
		"10000010",
		"10010000",
		"10011001",
		"10011100",
		"10100010",
		"10101001",
		"10101110",
		"10110011",
		"10110100",
		"10110111",
		"10110111",
		"10110101",
		"10110111",
		"10111001",
		"10111100",
		"10111110",
		"10111111",
		"11000000",
		"10111111",
		"10111101",
		"10100110",
		"01101100",
		"01000101",
		"01010010",
		"01111001",
		"10000100",
		"10000101",
		"10001111",
		"10011100",
		"10100011",
		"10101011",
		"10101111",
		"10101111",
		"10101111",
		"10101110",
		"10101110",
		"10101011",
		"10100010",
		"01110111",
		"10110011",
		"10101101",
		"10101110",
		"10101110",
		"10101111",
		"10110010",
		"10110100",
		"10110110",
		"10111000",
		"10111000",
		"10111010",
		"10110100",
		"10010010",
		"01011101",
		"01010010",
		"01010011",
		"01010011",
		"01010001",
		"01010011",
		"01010100",
		"01010100",
		"01010010",
		"01010010",
		"01010001",
		"01010000",
		"01010001",
		"01010011",
		"01010010",
		"01010001",
		"01010010",
		"01010011",
		"01010101",
		"01010011",
		"01011111",
		"01101100",
		"10010100",
		"10110101",
		"10101100",
		"01111001",
		"01010101",
		"01001011",
		"01001010",
		"01001111",
		"01010001",
		"01010010",
		"01010010",
		"01010001",
		"01010010",
		"01011010",
		"01101011",
		"01110010",
		"01100101",
		"01010101",
		"01010010",
		"01010110",
		"01011000",
		"01011000",
		"01011000",
		"01011000",
		"01011011",
		"01011100",
		"01011011",
		"01011101",
		"01011101",
		"01011101",
		"01100000",
		"01100001",
		"01100001",
		"01100001",
		"01100001",
		"01100001",
		"01100010",
		"01100011",
		"01100011",
		"01100011",
		"01100001",
		"01011111",
		"01011110",
		"01101110",
		"10011010",
		"11001010",
		"11011100",
		"11010100",
		"11001110",
		"11001010",
		"11000101",
		"11000001",
		"10110101",
		"10101010",
		"10010011",
		"01011000",
		"01011100",
		"01101110",
		"10000000",
		"10011110",
		"10100111",
		"11000101",
		"11000001",
		"10110111",
		"10010011",
		"10011101",
		"11001000",
		"10111100",
		"10110010",
		"10110001",
		"10111000",
		"10111011",
		"10111011",
		"10111011",
		"10110111",
		"10100001",
		"10001010",
		"10001100",
		"10010111",
		"10011110",
		"10100101",
		"10101001",
		"10101110",
		"10110001",
		"10110010",
		"10110100",
		"10110101",
		"10110111",
		"10111001",
		"10111001",
		"10111010",
		"10111101",
		"10111111",
		"11000000",
		"10111110",
		"10110110",
		"10011010",
		"01001110",
		"00101010",
		"01010110",
		"10000100",
		"10010001",
		"10001011",
		"10001101",
		"10011001",
		"10011101",
		"10100010",
		"10100010",
		"10100001",
		"10011110",
		"10011110",
		"10011110",
		"10100000",
		"10011111",
		"01111010",
		"10110111",
		"10110100",
		"10110101",
		"10110101",
		"10110111",
		"10110110",
		"10110110",
		"10110111",
		"10111001",
		"10111011",
		"10111011",
		"10111011",
		"10111010",
		"10001001",
		"01001010",
		"01000110",
		"01000111",
		"01011110",
		"10000011",
		"01111011",
		"01011101",
		"01010111",
		"01100000",
		"01011111",
		"01011000",
		"01001100",
		"01000010",
		"01000010",
		"01000011",
		"01001000",
		"01001001",
		"01010011",
		"01100110",
		"01010010",
		"01011010",
		"10010001",
		"10001110",
		"01011111",
		"01001110",
		"01010001",
		"01010011",
		"01011000",
		"01011001",
		"01011000",
		"01011010",
		"01011011",
		"01011001",
		"01010111",
		"01010111",
		"01010100",
		"01010010",
		"01010101",
		"01010101",
		"01010111",
		"01011010",
		"01011010",
		"01011011",
		"01011100",
		"01011011",
		"01011100",
		"01011100",
		"01011100",
		"01011101",
		"01011111",
		"01011111",
		"01100001",
		"01100001",
		"01100001",
		"01100000",
		"01100000",
		"01100001",
		"01100011",
		"01100010",
		"01100011",
		"01100010",
		"01100011",
		"01100010",
		"01100001",
		"01011111",
		"01011101",
		"01101000",
		"10001110",
		"10111101",
		"11001101",
		"11000011",
		"10111001",
		"10101100",
		"10010101",
		"10000110",
		"01110000",
		"01110011",
		"01001110",
		"01000001",
		"10001001",
		"10100110",
		"10001000",
		"10010101",
		"10011010",
		"10111000",
		"11000011",
		"10111111",
		"11001010",
		"10111001",
		"10110100",
		"10101000",
		"10110101",
		"11001001",
		"11001001",
		"11000100",
		"11000000",
		"10111010",
		"10101001",
		"10001011",
		"10010010",
		"10011110",
		"10100010",
		"10100011",
		"10100011",
		"10100101",
		"10101001",
		"10101011",
		"10101110",
		"10110011",
		"10110110",
		"10111000",
		"10111011",
		"10111100",
		"10111011",
		"10111010",
		"10110111",
		"10101000",
		"10000010",
		"00101100",
		"00011111",
		"01101110",
		"10010010",
		"10011001",
		"10010000",
		"10001000",
		"10001111",
		"10010110",
		"10010111",
		"10010110",
		"10010100",
		"10010011",
		"10010101",
		"10010100",
		"10010110",
		"10011011",
		"01111011",
		"10111100",
		"10111001",
		"10111011",
		"10111100",
		"10111110",
		"11000100",
		"11001010",
		"11001010",
		"11010001",
		"11001110",
		"11000101",
		"10111101",
		"10111100",
		"10011101",
		"01001110",
		"01000000",
		"01000111",
		"01110110",
		"10010101",
		"10010010",
		"10001010",
		"10001101",
		"10010101",
		"10011000",
		"10010110",
		"10001100",
		"01111001",
		"01100000",
		"01000111",
		"01000100",
		"01000101",
		"01010000",
		"01100101",
		"01010000",
		"01101111",
		"10000001",
		"01011011",
		"01010000",
		"01001111",
		"01010011",
		"01010110",
		"01010110",
		"01011000",
		"01011000",
		"01011000",
		"01011000",
		"01011000",
		"01010101",
		"01010011",
		"01010100",
		"01010101",
		"01010111",
		"01010110",
		"01010110",
		"01010111",
		"01011001",
		"01011010",
		"01011011",
		"01011001",
		"01011011",
		"01011100",
		"01011011",
		"01011100",
		"01011101",
		"01011110",
		"01011111",
		"01011110",
		"01011111",
		"01011111",
		"01100000",
		"01100000",
		"01100001",
		"01100001",
		"01100000",
		"01100000",
		"01011111",
		"01100001",
		"01011111",
		"01100001",
		"01100100",
		"01100000",
		"01011100",
		"01101000",
		"10001101",
		"10101000",
		"10001110",
		"01110011",
		"01011100",
		"01111011",
		"10000100",
		"10001000",
		"01110000",
		"01100001",
		"10010111",
		"10100110",
		"10010100",
		"10110000",
		"10100101",
		"10100110",
		"11000010",
		"11001001",
		"11001000",
		"11001111",
		"11001000",
		"10101111",
		"10111000",
		"11001110",
		"11010110",
		"11010100",
		"11001010",
		"10111111",
		"10111001",
		"10101011",
		"10001110",
		"10010100",
		"10011000",
		"10011101",
		"10100001",
		"10100110",
		"10101011",
		"10101111",
		"10110100",
		"10110101",
		"10110101",
		"10110111",
		"10111000",
		"10111001",
		"10111001",
		"10110010",
		"10101001",
		"10010111",
		"01100101",
		"00010110",
		"00110101",
		"10001100",
		"10011001",
		"10011011",
		"10010111",
		"10001011",
		"10000100",
		"10001010",
		"10001111",
		"10001111",
		"10001111",
		"10010011",
		"10010111",
		"10011101",
		"10100001",
		"10011111",
		"10000011",
		"10111111",
		"10111011",
		"10111110",
		"10111111",
		"11000000",
		"11000011",
		"11000101",
		"11000100",
		"11001011",
		"11001000",
		"10111100",
		"10110111",
		"10101110",
		"01110101",
		"00111111",
		"01000110",
		"01101111",
		"10001100",
		"10001100",
		"10001101",
		"10010111",
		"10011100",
		"10011111",
		"10100011",
		"10100100",
		"10100110",
		"10100111",
		"10011111",
		"10000011",
		"01000100",
		"00011100",
		"00011000",
		"00011100",
		"01100100",
		"10001100",
		"01100101",
		"01001110",
		"01010101",
		"01010001",
		"01010001",
		"01010100",
		"01010110",
		"01010111",
		"01011000",
		"01010111",
		"01010110",
		"01010100",
		"01010100",
		"01010101",
		"01010010",
		"01010100",
		"01010100",
		"01010010",
		"01010010",
		"01010011",
		"01010111",
		"01011000",
		"01011010",
		"01011010",
		"01011001",
		"01011010",
		"01011001",
		"01011011",
		"01011011",
		"01011011",
		"01011010",
		"01011011",
		"01011100",
		"01011101",
		"01100000",
		"01100001",
		"01100001",
		"01100010",
		"01100010",
		"01100001",
		"01100000",
		"01100000",
		"01011110",
		"01100000",
		"01100011",
		"01100100",
		"01100100",
		"01100010",
		"01100011",
		"01110000",
		"01010111",
		"00011101",
		"01100100",
		"10100001",
		"10001001",
		"10000011",
		"01110010",
		"01011010",
		"10000001",
		"10011101",
		"10000111",
		"10011101",
		"10101100",
		"10011010",
		"10010111",
		"11000000",
		"11001010",
		"11000000",
		"10111101",
		"10111110",
		"11000101",
		"11001111",
		"11010100",
		"11010010",
		"11001010",
		"11000011",
		"10111100",
		"10111000",
		"10011110",
		"10010100",
		"10011101",
		"10100011",
		"10100111",
		"10101100",
		"10110001",
		"10110110",
		"10111001",
		"10111000",
		"10111001",
		"10111001",
		"10111000",
		"10110110",
		"10110101",
		"10101100",
		"10100000",
		"10001000",
		"01000101",
		"00010000",
		"01011000",
		"10010101",
		"10011000",
		"10011001",
		"10011010",
		"10010111",
		"10010011",
		"10001101",
		"10001101",
		"10010000",
		"10010010",
		"10011001",
		"10011111",
		"10100111",
		"10101011",
		"10101000",
		"10000110",
		"11000001",
		"10111100",
		"10111011",
		"10111011",
		"10111001",
		"10111001",
		"11000011",
		"11001010",
		"11001110",
		"11010100",
		"11001001",
		"10111001",
		"10011001",
		"01000001",
		"00110000",
		"01110101",
		"10001101",
		"10001101",
		"10010010",
		"10011010",
		"10011101",
		"10100001",
		"10100100",
		"10100101",
		"10100101",
		"10100101",
		"10100110",
		"10101000",
		"10100110",
		"01110011",
		"00011000",
		"00010010",
		"00111000",
		"10001011",
		"10000000",
		"01011010",
		"01010010",
		"01010100",
		"01010100",
		"01010010",
		"01010100",
		"01010111",
		"01010110",
		"01010110",
		"01010110",
		"01010101",
		"01010100",
		"01010100",
		"01010011",
		"01010011",
		"01010100",
		"01010001",
		"01010011",
		"01011101",
		"01010100",
		"01010011",
		"01010110",
		"01010111",
		"01011010",
		"01011011",
		"01011001",
		"01011010",
		"01011010",
		"01011011",
		"01011011",
		"01011000",
		"01011000",
		"01011000",
		"01011001",
		"01011110",
		"01011111",
		"01100001",
		"01100000",
		"01100010",
		"01100001",
		"01100000",
		"01011111",
		"01011110",
		"01011111",
		"01100000",
		"01100001",
		"01100011",
		"01100001",
		"01100000",
		"01100001",
		"01100100",
		"01011011",
		"10000111",
		"10001101",
		"01110100",
		"01110001",
		"01101001",
		"01100000",
		"01101101",
		"01110111",
		"10001011",
		"10011101",
		"10101000",
		"10101110",
		"10101101",
		"10110111",
		"10111011",
		"11000000",
		"11001100",
		"11010100",
		"11010111",
		"11010100",
		"11001110",
		"11000101",
		"11000010",
		"11000100",
		"11000010",
		"10111010",
		"10110010",
		"10011111",
		"10100100",
		"10101000",
		"10101110",
		"10110011",
		"10110110",
		"10111000",
		"10111010",
		"10111010",
		"10111001",
		"10111000",
		"10110100",
		"10110000",
		"10101100",
		"10100100",
		"10001111",
		"01100100",
		"00100010",
		"00100011",
		"01111001",
		"10010110",
		"10010110",
		"10010110",
		"10011001",
		"10011011",
		"10100011",
		"10011110",
		"10010000",
		"10001101",
		"10010010",
		"10010110",
		"10011101",
		"10100011",
		"10101011",
		"10101000",
		"01111110",
		"11000000",
		"10111010",
		"10111010",
		"10111001",
		"10111001",
		"10111001",
		"11000000",
		"11001101",
		"11001101",
		"11001010",
		"11000011",
		"10101000",
		"01101001",
		"00111111",
		"01101000",
		"10001111",
		"10010000",
		"10010100",
		"10011010",
		"10011111",
		"10100010",
		"10100100",
		"10100011",
		"10100101",
		"10110000",
		"10110001",
		"10100101",
		"10100000",
		"10010010",
		"01100000",
		"00101111",
		"01000110",
		"10000101",
		"10010001",
		"01110011",
		"01010111",
		"01010001",
		"01010100",
		"01010001",
		"01010010",
		"01010101",
		"01010101",
		"01010101",
		"01010110",
		"01010110",
		"01010110",
		"01010100",
		"01010011",
		"01010100",
		"01010101",
		"01010011",
		"01011111",
		"01111011",
		"10001111",
		"10000111",
		"01101000",
		"01011001",
		"01011010",
		"01011001",
		"01011010",
		"01011011",
		"01011011",
		"01011100",
		"01011111",
		"01100010",
		"01100000",
		"01011100",
		"01010110",
		"01010101",
		"01010101",
		"01011001",
		"01011100",
		"01011101",
		"01011111",
		"01011111",
		"01100001",
		"01011110",
		"01011110",
		"01011111",
		"01011110",
		"01011101",
		"01011101",
		"01011011",
		"01011100",
		"01011100",
		"01011111",
		"01100100",
		"01100101",
		"01101010",
		"01101000",
		"01101001",
		"01100101",
		"01110111",
		"01110000",
		"10000000",
		"10011001",
		"10100101",
		"10101010",
		"10110000",
		"10111000",
		"10111101",
		"10111110",
		"11000110",
		"11010000",
		"11010110",
		"11010110",
		"11001111",
		"11000110",
		"11000001",
		"11000000",
		"11000010",
		"11000011",
		"10111111",
		"10111000",
		"10101010",
		"10100111",
		"10101001",
		"10101101",
		"10110011",
		"10111000",
		"10111010",
		"10111011",
		"10111011",
		"10111010",
		"10110110",
		"10101100",
		"10100110",
		"10011110",
		"10001111",
		"01100110",
		"00100110",
		"00001010",
		"00110011",
		"10000101",
		"10010101",
		"10010101",
		"10010100",
		"10010111",
		"10011000",
		"10011010",
		"10011010",
		"10010100",
		"10001010",
		"10001110",
		"10010111",
		"10011111",
		"10100101",
		"10101110",
		"10101011",
		"01111110",
		"10111111",
		"10111001",
		"10111001",
		"10111000",
		"10110110",
		"10110110",
		"10110111",
		"10110111",
		"10111000",
		"10110010",
		"10011001",
		"01100101",
		"01000101",
		"01101011",
		"10001011",
		"10001010",
		"10010000",
		"10011010",
		"10100000",
		"10100010",
		"10100010",
		"10100000",
		"10100110",
		"11000100",
		"11011011",
		"11010110",
		"10100111",
		"10001001",
		"01011011",
		"00011011",
		"00100110",
		"01110110",
		"10010111",
		"10000010",
		"01101001",
		"01010111",
		"01010011",
		"01010101",
		"01010010",
		"01010001",
		"01010001",
		"01010010",
		"01010101",
		"01010101",
		"01010100",
		"01010100",
		"01010001",
		"01010110",
		"01011001",
		"01010111",
		"01100010",
		"10001001",
		"10011011",
		"10111100",
		"10110100",
		"01110001",
		"01010111",
		"01011001",
		"01011000",
		"01010111",
		"01010111",
		"01011110",
		"01100010",
		"01100100",
		"01100101",
		"01100010",
		"01011110",
		"01011001",
		"01010111",
		"01010111",
		"01011000",
		"01011011",
		"01011110",
		"01011101",
		"01011100",
		"01011110",
		"01011111",
		"01100000",
		"01011110",
		"01011100",
		"01011100",
		"01011011",
		"01011001",
		"01011001",
		"01011001",
		"01011100",
		"01011100",
		"01011100",
		"01011101",
		"01100001",
		"01101001",
		"01111101",
		"10000010",
		"01111000",
		"10000000",
		"10010010",
		"10011111",
		"10100111",
		"10101100",
		"10110101",
		"10111010",
		"10111110",
		"11000100",
		"11000110",
		"11000111",
		"11000111",
		"11000010",
		"10111110",
		"10111101",
		"10111111",
		"11000001",
		"11000010",
		"11000011",
		"10111011",
		"10110010",
		"10101100",
		"10101111",
		"10110000",
		"10110010",
		"10110111",
		"10111001",
		"10111010",
		"10111010",
		"10111001",
		"10101111",
		"10100000",
		"10010110",
		"10000010",
		"01010111",
		"00100001",
		"00001010",
		"00001000",
		"01000100",
		"10001101",
		"10010110",
		"10010110",
		"10010100",
		"10010011",
		"10011000",
		"10011001",
		"10011011",
		"10010110",
		"10001001",
		"10001111",
		"10011010",
		"10100001",
		"10101000",
		"10101111",
		"10101100",
		"01100101",
		"10001100",
		"10000111",
		"10010010",
		"10011101",
		"10101011",
		"10110011",
		"10110011",
		"10110010",
		"10101001",
		"10000111",
		"01010110",
		"00111000",
		"01011001",
		"10000100",
		"10001001",
		"10001110",
		"10010110",
		"10011111",
		"10100001",
		"10011111",
		"10011101",
		"10100110",
		"11001001",
		"11100010",
		"11011101",
		"10110010",
		"01111100",
		"01001010",
		"00010100",
		"00010011",
		"01100110",
		"10010000",
		"10001110",
		"01110110",
		"01100001",
		"01010110",
		"01010100",
		"01010100",
		"01010011",
		"01010010",
		"01010001",
		"01010011",
		"01010100",
		"01010101",
		"01010010",
		"01001111",
		"01010101",
		"01011011",
		"01011010",
		"01011111",
		"10000100",
		"10011111",
		"11000000",
		"10111110",
		"10000100",
		"01010110",
		"01011000",
		"01011000",
		"01010111",
		"01010111",
		"01010100",
		"01011000",
		"01100000",
		"01100010",
		"01100000",
		"01011101",
		"01011010",
		"01011001",
		"01011001",
		"01011001",
		"01011001",
		"01011011",
		"01011101",
		"01011110",
		"01011101",
		"01011110",
		"01011110",
		"01100001",
		"01100001",
		"01100001",
		"01011111",
		"01011110",
		"01011101",
		"01011101",
		"01011011",
		"01011110",
		"01011101",
		"01011100",
		"01011101",
		"01011110",
		"01011111",
		"01011111",
		"01100100",
		"01101101",
		"01111000",
		"10001110",
		"10011101",
		"10100101",
		"10101011",
		"10110100",
		"10111001",
		"10111010",
		"10111010",
		"10111001",
		"10111001",
		"10111011",
		"10111110",
		"11000000",
		"10111111",
		"11000001",
		"11000001",
		"11000011",
		"11000100",
		"10111111",
		"10110101",
		"10101011",
		"10110011",
		"10110101",
		"10110101",
		"10110111",
		"10111010",
		"10111011",
		"10111000",
		"10110011",
		"10011011",
		"01111110",
		"01100010",
		"00110111",
		"00010001",
		"00000110",
		"00001001",
		"00000101",
		"01000101",
		"10001111",
		"10010110",
		"10010111",
		"10010101",
		"10010011",
		"10010100",
		"10011010",
		"10011100",
		"10011101",
		"10010101",
		"10010001",
		"10011011",
		"10100000",
		"10100011",
		"10101001",
		"10101001",
		"01011000",
		"01111101",
		"10000010",
		"10000101",
		"10001000",
		"10001101",
		"10011001",
		"10100101",
		"10100010",
		"01110100",
		"01000001",
		"00101001",
		"01001011",
		"10000010",
		"10000110",
		"10001001",
		"10010100",
		"10011110",
		"10100000",
		"10011101",
		"10100001",
		"10111110",
		"11010100",
		"11011101",
		"11000001",
		"10001010",
		"01010100",
		"00101100",
		"00001100",
		"00010010",
		"01011101",
		"01111011",
		"01100010",
		"01010100",
		"01011101",
		"01011101",
		"01010101",
		"01010100",
		"01010100",
		"01010100",
		"01010010",
		"01010000",
		"01010010",
		"01010001",
		"01010000",
		"01001111",
		"01010000",
		"01011010",
		"01011111",
		"01101011",
		"10000100",
		"10010101",
		"10111010",
		"11000001",
		"10001110",
		"01010111",
		"01010110",
		"01010110",
		"01011001",
		"01011011",
		"01011001",
		"01010111",
		"01010111",
		"01010101",
		"01011001",
		"01011110",
		"01011001",
		"01010111",
		"01010111",
		"01011000",
		"01011000",
		"01011000",
		"01011010",
		"01011100",
		"01011101",
		"01100000",
		"01100001",
		"01100001",
		"01100001",
		"01100010",
		"01100010",
		"01100010",
		"01100011",
		"01100101",
		"01100100",
		"01100000",
		"01011110",
		"01100000",
		"01011101",
		"01011110",
		"01011111",
		"01011111",
		"01011111",
		"01011110",
		"01011110",
		"01011100",
		"01100010",
		"01111011",
		"10011111",
		"10101101",
		"10101101",
		"10110010",
		"10110111",
		"10110100",
		"10110100",
		"10110100",
		"10110101",
		"10110111",
		"10111010",
		"10111101",
		"10111111",
		"10111110",
		"11000000",
		"11000010",
		"11000000",
		"10111000",
		"10110010",
		"10110011",
		"10110111",
		"10111001",
		"10111000",
		"10111010",
		"10111001",
		"10110111",
		"10101000",
		"01101010",
		"00110011",
		"00010111",
		"00001000",
		"00000101",
		"00000111",
		"00001000",
		"00000100",
		"00110010",
		"10001010",
		"10010110",
		"10010111",
		"10010101",
		"10010011",
		"10010000",
		"10010101",
		"10011010",
		"10011101",
		"10011100",
		"10011000",
		"10011011",
		"10100100",
		"10101001",
		"10101110",
		"10101011",
		"01100100",
		"10001101",
		"10010011",
		"10010110",
		"10010111",
		"10011010",
		"10011100",
		"10011111",
		"10100000",
		"10001001",
		"00111010",
		"00110110",
		"01111101",
		"10000110",
		"10001001",
		"10010010",
		"10011011",
		"10011100",
		"10010111",
		"10011000",
		"10100001",
		"10111001",
		"10111111",
		"10010100",
		"01011000",
		"00101110",
		"00010100",
		"00000111",
		"00100000",
		"01011101",
		"01100010",
		"01001001",
		"01001000",
		"01100000",
		"01011100",
		"01011010",
		"01010111",
		"01010100",
		"01010011",
		"01010011",
		"01010011",
		"01010001",
		"01010001",
		"01010001",
		"01010000",
		"01010000",
		"01010001",
		"01011101",
		"01101101",
		"01111001",
		"10001111",
		"10101101",
		"10111101",
		"10100000",
		"01011110",
		"01010100",
		"01010111",
		"01011001",
		"01011011",
		"01011011",
		"01011001",
		"01011011",
		"01011010",
		"01011000",
		"01011000",
		"01010111",
		"01011000",
		"01011000",
		"01010111",
		"01011000",
		"01011010",
		"01011001",
		"01011001",
		"01011100",
		"01011100",
		"01011101",
		"01100000",
		"01100011",
		"01100011",
		"01100010",
		"01100011",
		"01100100",
		"01100011",
		"01100101",
		"01100100",
		"01100110",
		"01100011",
		"01100011",
		"01011110",
		"01011101",
		"01100000",
		"01100000",
		"01011111",
		"01011111",
		"01011110",
		"01011110",
		"01011110",
		"01011011",
		"01100101",
		"10010100",
		"10101110",
		"10101100",
		"10101111",
		"10110001",
		"10110001",
		"10110100",
		"10110011",
		"10110100",
		"10110111",
		"10111011",
		"10111100",
		"10111010",
		"10111101",
		"10111111",
		"10111111",
		"10111010",
		"10110111",
		"10110100",
		"10110111",
		"10111010",
		"10111101",
		"10111011",
		"10111000",
		"10110101",
		"10010010",
		"00100100",
		"00000101",
		"00000111",
		"00000111",
		"00000111",
		"00001001",
		"00001001",
		"00000111",
		"00011110",
		"01111101",
		"10010100",
		"10010110",
		"10010101",
		"10010100",
		"10001110",
		"10000111",
		"10010010",
		"10011011",
		"10011101",
		"10011010",
		"10011010",
		"10100101",
		"10101101",
		"10110100",
		"10110010",
		"01101101",
		"10010101",
		"10010111",
		"10011100",
		"10011011",
		"10100000",
		"10100100",
		"10100110",
		"10101001",
		"10101000",
		"10001001",
		"01101000",
		"10000010",
		"10000101",
		"10001111",
		"10010110",
		"10010010",
		"10010101",
		"10011111",
		"10101010",
		"10100011",
		"10000010",
		"01011111",
		"00110100",
		"00010111",
		"00001100",
		"00000101",
		"00100100",
		"01100100",
		"01010110",
		"01001001",
		"01001000",
		"01100000",
		"01101101",
		"01100000",
		"01011001",
		"01010111",
		"01010101",
		"01010011",
		"01010011",
		"01010100",
		"01010001",
		"01010000",
		"01001101",
		"01001111",
		"01001110",
		"01001101",
		"01100001",
		"01111011",
		"01111101",
		"10100111",
		"10111010",
		"10101011",
		"01101110",
		"01010011",
		"01010101",
		"01011000",
		"01011001",
		"01011011",
		"01011110",
		"01011100",
		"01011101",
		"01100110",
		"01101000",
		"01011101",
		"01011000",
		"01011000",
		"01011001",
		"01011010",
		"01011010",
		"01011100",
		"01011100",
		"01011010",
		"01011001",
		"01011100",
		"01011011",
		"01011101",
		"01011111",
		"01100010",
		"01100011",
		"01100010",
		"01100100",
		"01100100",
		"01100011",
		"01100011",
		"01100100",
		"01100001",
		"01100010",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01100001",
		"01100000",
		"01100000",
		"01100000",
		"01011111",
		"01100001",
		"01100000",
		"01100000",
		"10000100",
		"10101111",
		"10101110",
		"10110001",
		"10110100",
		"10110101",
		"10110010",
		"10110011",
		"10110111",
		"10111011",
		"10111100",
		"10111001",
		"10111101",
		"11000000",
		"10111110",
		"10111101",
		"10111011",
		"10110111",
		"10110101",
		"10111101",
		"10111111",
		"10111110",
		"10111011",
		"10110010",
		"01100101",
		"00000101",
		"00000101",
		"00001000",
		"00001001",
		"00001010",
		"00001000",
		"00001000",
		"00000111",
		"00001100",
		"01011101",
		"10001100",
		"10010010",
		"10010101",
		"10010011",
		"10010011",
		"10001001",
		"10001000",
		"10010101",
		"10011011",
		"10011100",
		"10011011",
		"10100100",
		"10101101",
		"10110110",
		"10110100",
		"01101011",
		"10010100",
		"10010101",
		"10011011",
		"10011101",
		"10011111",
		"10100011",
		"10100111",
		"10101000",
		"10101000",
		"10100010",
		"01111100",
		"01111001",
		"10001000",
		"10001101",
		"10010110",
		"10110000",
		"11001101",
		"11000001",
		"10011010",
		"01110111",
		"01000010",
		"00011111",
		"00001110",
		"00001011",
		"00001000",
		"00110010",
		"01101110",
		"01011100",
		"01001111",
		"01001111",
		"01011100",
		"01101101",
		"01101110",
		"01011011",
		"01010111",
		"01010111",
		"01010100",
		"01010011",
		"01010010",
		"01010010",
		"01010001",
		"01001110",
		"01001110",
		"01001101",
		"01001100",
		"01011010",
		"01110101",
		"01110010",
		"10011100",
		"10110011",
		"10101110",
		"01110101",
		"01010101",
		"01010100",
		"01010101",
		"01010111",
		"01011000",
		"01011010",
		"01011101",
		"01011101",
		"01011110",
		"01100100",
		"01100001",
		"01011101",
		"01011101",
		"01011001",
		"01011011",
		"01011100",
		"01011011",
		"01011101",
		"01011101",
		"01011101",
		"01011101",
		"01011110",
		"01011101",
		"01011110",
		"01011101",
		"01100001",
		"01100010",
		"01100010",
		"01100100",
		"01100100",
		"01100011",
		"01100011",
		"01100100",
		"01100011",
		"01100010",
		"01100001",
		"01011111",
		"01011111",
		"01011110",
		"01100000",
		"01100001",
		"01100001",
		"01100010",
		"01100001",
		"01100011",
		"01100011",
		"01100000",
		"01100000",
		"10000011",
		"10101111",
		"10110000",
		"10110001",
		"10110010",
		"10101111",
		"10110010",
		"10110110",
		"10111000",
		"10111010",
		"10111011",
		"10111100",
		"10111111",
		"11000000",
		"11000001",
		"10111111",
		"10111101",
		"10110110",
		"10111100",
		"10111011",
		"10110111",
		"10110100",
		"10100110",
		"01000100",
		"00001010",
		"00000111",
		"00001000",
		"00001011",
		"00001110",
		"00010111",
		"00100101",
		"00110110",
		"01001010",
		"01101100",
		"10001000",
		"10001100",
		"10010000",
		"10010001",
		"10010000",
		"10001010",
		"01111010",
		"10000000",
		"10010111",
		"10011010",
		"10011001",
		"10100100",
		"10101111",
		"10110111",
		"10110011",
		"01100010",
		"10001100",
		"10010000",
		"10011000",
		"10011010",
		"10011100",
		"10100001",
		"10100110",
		"10101001",
		"10100101",
		"10100010",
		"10000011",
		"01111001",
		"10001100",
		"10101110",
		"11010011",
		"11010110",
		"10110000",
		"01110110",
		"01001001",
		"00100010",
		"00010001",
		"00001011",
		"00001010",
		"00000110",
		"00101000",
		"10000110",
		"01101110",
		"01011100",
		"01010101",
		"01010111",
		"01100000",
		"01011110",
		"01011010",
		"01010110",
		"01010111",
		"01010110",
		"01010101",
		"01010101",
		"01010100",
		"01010011",
		"01010010",
		"01010000",
		"01001111",
		"01001110",
		"01010100",
		"01111101",
		"01111001",
		"10001011",
		"10101100",
		"10110010",
		"10000000",
		"01011001",
		"01010110",
		"01010101",
		"01010101",
		"01010110",
		"01010110",
		"01011001",
		"01011011",
		"01011101",
		"01011110",
		"01011111",
		"01100000",
		"01100000",
		"01011111",
		"01011011",
		"01011010",
		"01011100",
		"01011101",
		"01011110",
		"01011111",
		"01011111",
		"01100000",
		"01100010",
		"01011111",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01100010",
		"01100011",
		"01100100",
		"01100100",
		"01100101",
		"01100101",
		"01100100",
		"01100011",
		"01100010",
		"01100001",
		"01100001",
		"01100001",
		"01100001",
		"01100010",
		"01100000",
		"01100001",
		"01100001",
		"01100010",
		"01100011",
		"01100011",
		"01100101",
		"01100100",
		"10001000",
		"10100100",
		"10101110",
		"10101100",
		"10101101",
		"10101110",
		"10110001",
		"10110110",
		"10111001",
		"10111011",
		"10111111",
		"11000011",
		"11000001",
		"10111101",
		"10110100",
		"10101000",
		"10000111",
		"01100010",
		"01101101",
		"01110111",
		"01111101",
		"10000100",
		"10000100",
		"10000001",
		"01100100",
		"01000011",
		"00111000",
		"00110111",
		"01011010",
		"01111010",
		"10000110",
		"10010010",
		"10010011",
		"10010100",
		"10010110",
		"10010101",
		"10010111",
		"10010111",
		"10010011",
		"10000111",
		"01111111",
		"10001111",
		"10011000",
		"10011000",
		"10100011",
		"10101101",
		"10110111",
		"10110101",
		"01100010",
		"10001001",
		"10001110",
		"10010100",
		"10011001",
		"10011010",
		"10100001",
		"10100100",
		"10100110",
		"10011111",
		"10011101",
		"10001000",
		"10000010",
		"10011101",
		"10111110",
		"10110011",
		"10000111",
		"01010011",
		"00101100",
		"00010011",
		"00001101",
		"00001011",
		"00001010",
		"00000100",
		"00010100",
		"01100010",
		"10000011",
		"01101001",
		"01011011",
		"01010101",
		"01010010",
		"01010100",
		"01010010",
		"01001111",
		"01010011",
		"01010011",
		"01010100",
		"01010011",
		"01010100",
		"01010100",
		"01010010",
		"01001111",
		"01001111",
		"01001101",
		"01001011",
		"01110011",
		"10001000",
		"10010011",
		"10101100",
		"10111010",
		"10011100",
		"01100000",
		"01011010",
		"01011000",
		"01011000",
		"01010111",
		"01010110",
		"01010110",
		"01011001",
		"01011100",
		"01011101",
		"01011111",
		"01100000",
		"01100010",
		"01100001",
		"01011111",
		"01011110",
		"01011000",
		"01011010",
		"01011101",
		"01011101",
		"01011110",
		"01100000",
		"01100000",
		"01100001",
		"01100011",
		"01100010",
		"01100010",
		"01100001",
		"01100010",
		"01100010",
		"01100010",
		"01100100",
		"01100101",
		"01100111",
		"01100110",
		"01100101",
		"01100101",
		"01100100",
		"01100001",
		"01100011",
		"01100010",
		"01100010",
		"01100010",
		"01100010",
		"01100000",
		"01100001",
		"01100011",
		"01101010",
		"01101100",
		"01100101",
		"01100100",
		"01101000",
		"01110011",
		"10001000",
		"10100111",
		"10100111",
		"10101010",
		"10101101",
		"10110100",
		"10111100",
		"11000000",
		"10111000",
		"10101001",
		"10010111",
		"10000111",
		"01111001",
		"01110011",
		"01100001",
		"01011011",
		"01100111",
		"01110101",
		"10000001",
		"10001000",
		"10010100",
		"10011100",
		"10100001",
		"10100100",
		"10010111",
		"10000011",
		"01111001",
		"10000001",
		"10001111",
		"10011000",
		"10011011",
		"10011001",
		"10011100",
		"10100000",
		"10100000",
		"10100000",
		"10100001",
		"10011101",
		"10010101",
		"10001111",
		"10010011",
		"10011000",
		"10100010",
		"10101001",
		"10110010",
		"10110010",
		"01101010",
		"10001111",
		"10001010",
		"10010011",
		"10010110",
		"10011001",
		"10100001",
		"10100010",
		"10011111",
		"10011010",
		"10001001",
		"01001000",
		"01001111",
		"01111011",
		"01111111",
		"01100010",
		"00111000",
		"00011001",
		"00001111",
		"00001100",
		"00001011",
		"00001000",
		"00000100",
		"00111100",
		"01111000",
		"01101100",
		"01110000",
		"01100000",
		"01010101",
		"01010010",
		"01010000",
		"01001111",
		"01001110",
		"01001100",
		"01001110",
		"01010001",
		"01010011",
		"01010010",
		"01010100",
		"01010011",
		"01010010",
		"01010000",
		"01001110",
		"01001011",
		"01011110",
		"10000100",
		"10001001",
		"10100111",
		"10111110",
		"10111010",
		"10000001",
		"01011100",
		"01011111",
		"01011001",
		"01011000",
		"01011001",
		"01011000",
		"01011000",
		"01011001",
		"01011011",
		"01011100",
		"01011100",
		"01011110",
		"01100000",
		"01100011",
		"01100110",
		"01100110",
		"01011101",
		"01011000",
		"01011101",
		"01011100",
		"01011110",
		"01100001",
		"01100000",
		"01100001",
		"01100001",
		"01100001",
		"01100010",
		"01100011",
		"01100010",
		"01100000",
		"01100001",
		"01100010",
		"01100100",
		"01100101",
		"01100011",
		"01100101",
		"01100111",
		"01100101",
		"01100100",
		"01100011",
		"01100011",
		"01100100",
		"01100010",
		"01100000",
		"01100010",
		"01100000",
		"01100001",
		"01100011",
		"01100101",
		"01100101",
		"01100110",
		"01100110",
		"01101011",
		"01011101",
		"01110101",
		"10011111",
		"10100011",
		"10101001",
		"10110010",
		"10101001",
		"10010010",
		"01110110",
		"01101010",
		"01101000",
		"01101010",
		"01110010",
		"01110001",
		"01110010",
		"01110100",
		"01111011",
		"10000110",
		"10010010",
		"10010111",
		"10011011",
		"10011101",
		"10100000",
		"10100001",
		"10100110",
		"10100110",
		"10100001",
		"10010101",
		"10010000",
		"10011000",
		"10011011",
		"10011110",
		"10100101",
		"10100111",
		"10101001",
		"10101000",
		"10101000",
		"10100011",
		"10011111",
		"10011101",
		"10011000",
		"10010011",
		"10011001",
		"10100000",
		"10100110",
		"10101000",
		"01101011",
		"10001101",
		"10001001",
		"10010011",
		"10010101",
		"10011001",
		"10011011",
		"10011010",
		"10010111",
		"10010001",
		"01011001",
		"00010010",
		"00001101",
		"00011010",
		"00100001",
		"00011000",
		"00001101",
		"00001011",
		"00001011",
		"00001101",
		"00001001",
		"00010001",
		"01100000",
		"10101101",
		"10000011",
		"01011001",
		"01100000",
		"01010111",
		"01010010",
		"01010000",
		"01010000",
		"01001111",
		"01010001",
		"01001111",
		"01001110",
		"01010000",
		"01010011",
		"01010001",
		"01010001",
		"01010001",
		"01010001",
		"01010000",
		"01001111",
		"01010001",
		"10000000",
		"10000111",
		"10011001",
		"10101111",
		"10111010",
		"10110001",
		"01101011",
		"01011101",
		"01100001",
		"01011011",
		"01011000",
		"01011000",
		"01011000",
		"01011000",
		"01011000",
		"01011011",
		"01011101",
		"01011110",
		"01100001",
		"01100100",
		"01110011",
		"10000000",
		"10001010",
		"01111100",
		"01011100",
		"01011000",
		"01011011",
		"01011101",
		"01011111",
		"01100000",
		"01011111",
		"01011111",
		"01100000",
		"01100001",
		"01100011",
		"01100010",
		"01100000",
		"01100000",
		"01100000",
		"01100100",
		"01100010",
		"01100011",
		"01100101",
		"01100101",
		"01100101",
		"01100110",
		"01100100",
		"01100010",
		"01100100",
		"01100010",
		"01100010",
		"01100001",
		"01100011",
		"01100011",
		"01100100",
		"01100100",
		"01100101",
		"01100111",
		"01101001",
		"01100110",
		"01011110",
		"01011100",
		"01101100",
		"10010100",
		"10001011",
		"01110010",
		"01010110",
		"01000100",
		"01000001",
		"01000010",
		"01010101",
		"01101111",
		"01111010",
		"01110001",
		"01101101",
		"01110101",
		"10000110",
		"10010011",
		"10011001",
		"10011011",
		"10011111",
		"10100001",
		"10100010",
		"10100011",
		"10101010",
		"10100111",
		"10100111",
		"10100111",
		"10011111",
		"10011001",
		"10011110",
		"10100110",
		"10101101",
		"10110010",
		"10110100",
		"10110100",
		"10110000",
		"10101000",
		"10100101",
		"10100101",
		"10100010",
		"10011110",
		"10011100",
		"10011001",
		"10011101",
		"10100001",
		"01100011",
		"10001011",
		"10001100",
		"10010001",
		"10010101",
		"10011001",
		"10010101",
		"10001101",
		"10000101",
		"01101001",
		"00100110",
		"00010010",
		"00010000",
		"00001011",
		"00001010",
		"00001010",
		"00001100",
		"00001101",
		"00001111",
		"00001110",
		"00011100",
		"01111011",
		"10111000",
		"10101111",
		"01101110",
		"01010100",
		"01010011",
		"01010010",
		"01010010",
		"01010010",
		"01010001",
		"01010001",
		"01001111",
		"01010001",
		"01010001",
		"01010000",
		"01001111",
		"01010000",
		"01010000",
		"01010000",
		"01010000",
		"01001111",
		"01001111",
		"01110010",
		"01111101",
		"10001101",
		"10100110",
		"10111110",
		"10111101",
		"10100010",
		"01100000",
		"01100011",
		"01100010",
		"01011100",
		"01011001",
		"01011000",
		"01011011",
		"01011011",
		"01011011",
		"01011011",
		"01011111",
		"01100001",
		"01100000",
		"01100111",
		"01110010",
		"01111000",
		"10000111",
		"10011100",
		"01110110",
		"01010111",
		"01011010",
		"01011010",
		"01011100",
		"01011101",
		"01100000",
		"01011110",
		"01011101",
		"01011111",
		"01100010",
		"01100000",
		"01100000",
		"01011110",
		"01011110",
		"01100010",
		"01100110",
		"01100010",
		"01100010",
		"01100011",
		"01100101",
		"01100110",
		"01101000",
		"01100110",
		"01100011",
		"01100001",
		"01100010",
		"01100100",
		"01100111",
		"01101011",
		"01100110",
		"01100110",
		"01100101",
		"01100111",
		"01100111",
		"01100001",
		"01011111",
		"01011111",
		"01011101",
		"01100110",
		"01010000",
		"00011001",
		"00011011",
		"00101001",
		"00111100",
		"01001000",
		"01010100",
		"01011110",
		"01011001",
		"01100011",
		"01110011",
		"01111111",
		"10001001",
		"10010000",
		"10011000",
		"10011001",
		"10011101",
		"10100001",
		"10100100",
		"10101000",
		"10101010",
		"10101011",
		"10101100",
		"10101011",
		"10101000",
		"10100101",
		"10101001",
		"10110001",
		"10111011",
		"11000011",
		"11001000",
		"11000111",
		"10111111",
		"10110111",
		"10101100",
		"10101001",
		"10101000",
		"10100011",
		"10100111",
		"10100010",
		"10011111",
		"10011101",
		"01011110",
		"10000111",
		"10001011",
		"10001100",
		"10110010",
		"10111000",
		"10000101",
		"01101101",
		"01010000",
		"00100001",
		"00010011",
		"00010011",
		"00010010",
		"00010001",
		"00010100",
		"00010111",
		"00011001",
		"00011010",
		"00011000",
		"00011111",
		"01110010",
		"10101111",
		"10101010",
		"10011010",
		"01100110",
		"01001110",
		"01001111",
		"01010001",
		"01010011",
		"01010011",
		"01010010",
		"01010001",
		"01010000",
		"01001111",
		"01001111",
		"01001111",
		"01010000",
		"01010001",
		"01001111",
		"01010001",
		"01001111",
		"01010000",
		"01100101",
		"10001000",
		"10001110",
		"10011001",
		"10110001",
		"11000100",
		"11000101",
		"10100101",
		"01100001",
		"01100011",
		"01100110",
		"01100001",
		"01011011",
		"01011010",
		"01011011",
		"01011110",
		"01011111",
		"01011100",
		"01011111",
		"01100010",
		"01100100",
		"01100100",
		"01100101",
		"01100001",
		"01100111",
		"10000000",
		"10010001",
		"01100111",
		"01010100",
		"01011001",
		"01011011",
		"01011101",
		"01011101",
		"01011110",
		"01011110",
		"01100000",
		"01100010",
		"01100011",
		"01100010",
		"01100001",
		"01011111",
		"01100001",
		"01101000",
		"01100001",
		"01100010",
		"01100101",
		"01101011",
		"01110001",
		"01101001",
		"01100100",
		"01100011",
		"01100100",
		"01101110",
		"01111001",
		"01110110",
		"01111010",
		"10000111",
		"01110111",
		"01101000",
		"01100101",
		"01100100",
		"01101010",
		"01100111",
		"01100001",
		"01011110",
		"01011110",
		"01100000",
		"00101111",
		"00001110",
		"00100000",
		"00111001",
		"01001111",
		"01011101",
		"01010110",
		"01010011",
		"01100111",
		"01110010",
		"10000001",
		"10001100",
		"10001111",
		"10010110",
		"10011010",
		"10011101",
		"10100001",
		"10100111",
		"10101010",
		"10101010",
		"10101100",
		"10101111",
		"10110001",
		"10101110",
		"10101010",
		"10101110",
		"10110101",
		"10110111",
		"10111000",
		"10111010",
		"10111101",
		"11000111",
		"11000000",
		"10110111",
		"10111011",
		"10111111",
		"10111010",
		"10101100",
		"10100101",
		"10100100",
		"10100001",
		"01101101",
		"10011011",
		"10010111",
		"10011111",
		"11000110",
		"10110111",
		"10010011",
		"10001010",
		"01111011",
		"01101000",
		"01100011",
		"01010101",
		"01000000",
		"00100100",
		"00010111",
		"00011010",
		"00011111",
		"00011111",
		"00011111",
		"01101000",
		"10101101",
		"10101011",
		"10011110",
		"10010100",
		"01110110",
		"01001110",
		"01010001",
		"01010001",
		"01010010",
		"01010010",
		"01010010",
		"01010000",
		"01001111",
		"01001110",
		"01010000",
		"01010000",
		"01010001",
		"01010001",
		"01001111",
		"01010010",
		"01010110",
		"01111010",
		"10001011",
		"01111110",
		"10011000",
		"10011100",
		"10111010",
		"11000111",
		"11001010",
		"10111110",
		"01111100",
		"01011111",
		"01100001",
		"01011101",
		"01011100",
		"01011010",
		"01011010",
		"01011110",
		"01011100",
		"01011100",
		"01011111",
		"01100001",
		"01100001",
		"01100011",
		"01100111",
		"01100011",
		"01100000",
		"01100001",
		"01101100",
		"10010000",
		"01100101",
		"01011000",
		"01011010",
		"01011011",
		"01011100",
		"01011111",
		"01100000",
		"01100010",
		"01100000",
		"01100011",
		"01100001",
		"01100010",
		"01100010",
		"01100000",
		"01100000",
		"01100010",
		"01100100",
		"01100110",
		"01111110",
		"10101100",
		"10101011",
		"10011100",
		"01111011",
		"01101100",
		"10001011",
		"10010101",
		"10011101",
		"10101011",
		"10101100",
		"10011000",
		"01101111",
		"01100100",
		"01100100",
		"10010011",
		"10000110",
		"01100101",
		"01011110",
		"01011110",
		"01100010",
		"01100001",
		"00100001",
		"00010001",
		"00100001",
		"00111011",
		"01000100",
		"01001000",
		"01010101",
		"01100100",
		"01110001",
		"01111101",
		"10001000",
		"10001111",
		"10010110",
		"10011010",
		"10011111",
		"10100101",
		"10100111",
		"10101000",
		"10101110",
		"10110001",
		"10110100",
		"10110110",
		"10110010",
		"10101100",
		"10101011",
		"10111100",
		"10111001",
		"10110010",
		"10101011",
		"10100110",
		"10101010",
		"10101001",
		"10111001",
		"11001110",
		"11010101",
		"11011000",
		"11001000",
		"10101111",
		"10100110",
		"10100101",
		"10001011",
		"11000011",
		"10111100",
		"10111010",
		"10111000",
		"10111001",
		"10111011",
		"10111011",
		"10111100",
		"10111010",
		"10110111",
		"10101110",
		"10100001",
		"10000101",
		"01001111",
		"00101000",
		"00011111",
		"00011011",
		"01001110",
		"10100100",
		"10101100",
		"10100100",
		"10010111",
		"10010001",
		"10001101",
		"01010001",
		"01001111",
		"01010100",
		"01010010",
		"01010000",
		"01010000",
		"01001111",
		"01001111",
		"01001101",
		"01001101",
		"01001110",
		"01010000",
		"01010000",
		"01010010",
		"01000111",
		"01101101",
		"10001100",
		"10000101",
		"10010000",
		"10100100",
		"10100011",
		"10110011",
		"11001000",
		"11001110",
		"11000111",
		"10100000",
		"01011011",
		"01011001",
		"01011001",
		"01011001",
		"01011000",
		"01011001",
		"01011011",
		"01011011",
		"01011100",
		"01011111",
		"01100000",
		"01011110",
		"01100011",
		"01100111",
		"01100101",
		"01100010",
		"01100001",
		"01011110",
		"01110001",
		"10001011",
		"01010110",
		"01011000",
		"01011011",
		"01011101",
		"01011101",
		"01011110",
		"01100001",
		"01100010",
		"01100010",
		"01100100",
		"01100100",
		"01100010",
		"01100001",
		"01100011",
		"01100101",
		"01100110",
		"01100100",
		"10000001",
		"11000111",
		"11010100",
		"11010010",
		"11000010",
		"10100001",
		"10101100",
		"11000100",
		"11001001",
		"11001100",
		"10111101",
		"10011110",
		"01110100",
		"01100100",
		"01101000",
		"10100111",
		"10011111",
		"10000001",
		"01101010",
		"01100000",
		"01100000",
		"01101001",
		"01010000",
		"00010000",
		"00010111",
		"00100000",
		"00101010",
		"00111100",
		"01011000",
		"01101110",
		"01110110",
		"01111101",
		"10001001",
		"10001111",
		"10010100",
		"10011001",
		"10100001",
		"10100011",
		"10100110",
		"10101011",
		"10110101",
		"10111111",
		"11000001",
		"10110110",
		"10110000",
		"10101100",
		"10100111",
		"10111100",
		"11001000",
		"10110110",
		"10100100",
		"10011101",
		"10010110",
		"10011100",
		"10110001",
		"11001110",
		"11011101",
		"11100000",
		"11010101",
		"10111000",
		"10101111",
		"10101011",
		"10001011",
		"11000100",
		"10111111",
		"10111110",
		"10111100",
		"10111100",
		"10111100",
		"10111011",
		"10111011",
		"10111010",
		"10111000",
		"10101110",
		"10011101",
		"10001110",
		"01110100",
		"01010000",
		"00110011",
		"00101100",
		"10001011",
		"10101100",
		"10100011",
		"10011111",
		"10010101",
		"10001111",
		"10010101",
		"01101010",
		"01000101",
		"01010000",
		"01010011",
		"01010000",
		"01010001",
		"01001110",
		"01001100",
		"01001011",
		"01010011",
		"01010011",
		"01000100",
		"01001111",
		"01011110",
		"00110100",
		"01110100",
		"01111111",
		"01100110",
		"10010001",
		"10100000",
		"10100001",
		"10101100",
		"11000001",
		"11001000",
		"10111001",
		"10101100",
		"10000101",
		"01101101",
		"01011000",
		"01010101",
		"01010110",
		"01011000",
		"01011011",
		"01011100",
		"01011011",
		"01011100",
		"01011110",
		"01100001",
		"01100011",
		"01100110",
		"01101101",
		"01101100",
		"01101100",
		"01100100",
		"01011110",
		"10000100",
		"01110011",
		"01010110",
		"01011000",
		"01011011",
		"01011011",
		"01011101",
		"01011111",
		"01100000",
		"01100011",
		"01100101",
		"01100011",
		"01100011",
		"01100011",
		"01100010",
		"01100100",
		"01101010",
		"01100111",
		"01111011",
		"11000010",
		"11010110",
		"11010110",
		"11010101",
		"11001001",
		"11000100",
		"11010011",
		"11011001",
		"11011001",
		"11010110",
		"10101110",
		"01110000",
		"01100110",
		"01111011",
		"10101110",
		"10011001",
		"10001110",
		"01110110",
		"01100111",
		"01100001",
		"01100100",
		"01101001",
		"00101110",
		"00001111",
		"00011010",
		"00100111",
		"00111010",
		"01010000",
		"01101110",
		"01111100",
		"10000011",
		"10001010",
		"10010000",
		"10010111",
		"10011000",
		"10100000",
		"10100010",
		"10100111",
		"10110010",
		"11000000",
		"11001001",
		"11001010",
		"11000000",
		"10110011",
		"10101011",
		"10101000",
		"10110100",
		"10110101",
		"11000011",
		"10101100",
		"10010010",
		"10010010",
		"10011110",
		"10110000",
		"11001000",
		"11010111",
		"11010011",
		"10111000",
		"10011000",
		"10001010",
		"10001100",
		"10000111",
		"11000101",
		"10111111",
		"11000000",
		"10111110",
		"10111110",
		"10111101",
		"10111100",
		"10111010",
		"10111001",
		"10110011",
		"10100111",
		"10010010",
		"01111010",
		"01100000",
		"01001011",
		"00110011",
		"01011001",
		"10101000",
		"10100111",
		"10011110",
		"10010101",
		"10010001",
		"10001001",
		"10001111",
		"10011100",
		"01010110",
		"01000111",
		"01010011",
		"01010000",
		"01010001",
		"01001100",
		"01010001",
		"01111011",
		"01110001",
		"01101000",
		"01110111",
		"01111000",
		"01111010",
		"01111010",
		"01111110",
		"10000101",
		"01110011",
		"10000100",
		"01111010",
		"10001010",
		"10101010",
		"10110110",
		"10110011",
		"10011100",
		"10101000",
		"10110111",
		"10100010",
		"01111000",
		"01010110",
		"01010001",
		"01010110",
		"01011010",
		"01011100",
		"01011101",
		"01011100",
		"01011101",
		"01011111",
		"01100001",
		"01100011",
		"01101111",
		"10000010",
		"10001001",
		"01101101",
		"01100000",
		"01100101",
		"01111111",
		"01010101",
		"01010110",
		"01011001",
		"01011010",
		"01011100",
		"01011101",
		"01100001",
		"01100010",
		"01100101",
		"01100100",
		"01100001",
		"01100010",
		"01100010",
		"01100100",
		"01101001",
		"01101100",
		"10001010",
		"10111001",
		"11001100",
		"11011010",
		"11010110",
		"11001011",
		"11000010",
		"11000101",
		"11010011",
		"11010100",
		"11001101",
		"10100000",
		"01101100",
		"01110010",
		"01111001",
		"01111111",
		"01111000",
		"01110101",
		"01101101",
		"01100110",
		"01100000",
		"01100011",
		"01101001",
		"01001110",
		"00010001",
		"00011001",
		"00100101",
		"00111100",
		"01001101",
		"01100101",
		"01111101",
		"10001000",
		"10001110",
		"10010001",
		"10010100",
		"10011010",
		"10011110",
		"10100011",
		"10101001",
		"10110110",
		"11001000",
		"11001111",
		"11010000",
		"11001100",
		"10110110",
		"10101001",
		"10101000",
		"10110000",
		"10100110",
		"10100011",
		"10110111",
		"10100111",
		"10011100",
		"10011110",
		"10100110",
		"10100000",
		"10000010",
		"01100101",
		"01101000",
		"01110110",
		"10000100",
		"10010110",
		"10000111",
		"11001000",
		"11000001",
		"11000001",
		"11000001",
		"10111111",
		"10111101",
		"10111100",
		"10111010",
		"10110101",
		"10101011",
		"10011010",
		"10000001",
		"01100101",
		"01001011",
		"00111000",
		"00100011",
		"01110010",
		"10101100",
		"10100100",
		"10011011",
		"10010011",
		"10001100",
		"10000000",
		"10010000",
		"10100111",
		"10001111",
		"01000110",
		"01001011",
		"01010000",
		"01001100",
		"01011001",
		"10010111",
		"10101011",
		"10011001",
		"01111111",
		"01111110",
		"10001100",
		"10010110",
		"10010100",
		"10001001",
		"10000011",
		"10011011",
		"10011110",
		"01111011",
		"10001000",
		"10110000",
		"10101101",
		"10101001",
		"10101101",
		"10101010",
		"10111010",
		"10101001",
		"10100000",
		"10100001",
		"01110010",
		"01001111",
		"01010110",
		"01011100",
		"01011100",
		"01011101",
		"01011111",
		"01100000",
		"01100001",
		"01100110",
		"01101110",
		"01111011",
		"10010000",
		"10000000",
		"01100111",
		"01011101",
		"01101010",
		"01100010",
		"01010101",
		"01011000",
		"01011010",
		"01011100",
		"01011110",
		"01100000",
		"01100011",
		"01100011",
		"01100010",
		"01100011",
		"01100011",
		"01100011",
		"01100011",
		"01101001",
		"01111010",
		"10010011",
		"10110111",
		"11000101",
		"11010110",
		"11011001",
		"11000000",
		"10100110",
		"10110100",
		"11001110",
		"11001110",
		"10110101",
		"10000000",
		"01101011",
		"01110111",
		"01100111",
		"01011110",
		"01100011",
		"01101000",
		"01101100",
		"01100011",
		"01100001",
		"01100010",
		"01101010",
		"01100101",
		"00100001",
		"00010100",
		"00101000",
		"00111100",
		"01001011",
		"01011010",
		"01111010",
		"10000111",
		"10001101",
		"10010000",
		"10010101",
		"10011101",
		"10011111",
		"10100100",
		"10101010",
		"10111100",
		"11001111",
		"11010101",
		"11010100",
		"11001110",
		"10111010",
		"10100111",
		"10100101",
		"10100111",
		"10110001",
		"10100110",
		"10011001",
		"10101111",
		"11001000",
		"10100110",
		"01110111",
		"01011101",
		"01011000",
		"01110000",
		"10000110",
		"10010010",
		"10010111",
		"10011100",
		"10001001",
		"11001001",
		"11000011",
		"11000001",
		"11000010",
		"11000001",
		"10111110",
		"10111101",
		"10111011",
		"10110011",
		"10100011",
		"10000111",
		"01100011",
		"01000110",
		"00101001",
		"00010110",
		"00010111",
		"10000110",
		"10101110",
		"10100010",
		"10011100",
		"10010000",
		"10000000",
		"01111101",
		"10010100",
		"10100011",
		"10101110",
		"01110110",
		"00111111",
		"01001011",
		"01011101",
		"10011110",
		"10101110",
		"10011100",
		"10001010",
		"10000101",
		"01111111",
		"10001001",
		"10010100",
		"10010111",
		"10010000",
		"10000101",
		"10001101",
		"10011111",
		"10001100",
		"10010000",
		"10111111",
		"10111000",
		"10110101",
		"11001000",
		"11000100",
		"10110111",
		"10110101",
		"10110101",
		"10110010",
		"10110110",
		"01110011",
		"01001111",
		"01011000",
		"01011001",
		"01011110",
		"01011110",
		"01100000",
		"01100001",
		"01100110",
		"01111000",
		"10010000",
		"10100010",
		"10010001",
		"01101110",
		"01100011",
		"01011110",
		"01101001",
		"01010110",
		"01010111",
		"01011001",
		"01011100",
		"01011110",
		"01100000",
		"01100001",
		"01100010",
		"01100010",
		"01100010",
		"01100010",
		"01100011",
		"01100101",
		"01101010",
		"10000000",
		"10010110",
		"10110001",
		"11000001",
		"11001110",
		"11000000",
		"10011101",
		"10001010",
		"10101111",
		"10111010",
		"10101011",
		"10001011",
		"01101110",
		"01110001",
		"01110011",
		"01100010",
		"01011110",
		"01100001",
		"01100010",
		"01100001",
		"01100010",
		"01100000",
		"01100010",
		"01101111",
		"01110011",
		"00110100",
		"00010010",
		"00101000",
		"00111100",
		"01000111",
		"01011100",
		"01111100",
		"10001000",
		"10001101",
		"10010001",
		"10011000",
		"10011110",
		"10100010",
		"10100001",
		"10101011",
		"11000100",
		"11010011",
		"11011001",
		"11011000",
		"11010100",
		"10111001",
		"10100101",
		"10100101",
		"10100101",
		"10101001",
		"10011111",
		"10000111",
		"01110111",
		"01111100",
		"01100101",
		"01011001",
		"01100010",
		"01110101",
		"10001101",
		"10010110",
		"10010110",
		"10011110",
		"10100000",
		"10001000",
		"11000111",
		"11000010",
		"11000001",
		"11000000",
		"11000000",
		"10111111",
		"10111011",
		"10110110",
		"10101000",
		"10000101",
		"01011001",
		"00110110",
		"00011100",
		"00010000",
		"00001010",
		"00100110",
		"10011010",
		"10101100",
		"10100010",
		"10011100",
		"10010010",
		"10001001",
		"10010110",
		"10011111",
		"10100101",
		"10101001",
		"10101011",
		"01011110",
		"01001100",
		"10010011",
		"10101001",
		"10011110",
		"10001011",
		"10000010",
		"10000111",
		"10001100",
		"10010101",
		"10011101",
		"10100000",
		"10100011",
		"10100010",
		"10011111",
		"10100001",
		"10011011",
		"10011011",
		"10110011",
		"10110010",
		"10110100",
		"10110010",
		"10110010",
		"10110101",
		"10111000",
		"10110111",
		"10101101",
		"10110111",
		"10101111",
		"01011111",
		"01010110",
		"01011010",
		"01011110",
		"01100000",
		"01100001",
		"01100011",
		"01101001",
		"10000010",
		"10111100",
		"11001101",
		"10111110",
		"10001100",
		"01101001",
		"01011111",
		"01100100",
		"01011001",
		"01010101",
		"01011001",
		"01011000",
		"01011100",
		"01011110",
		"01011111",
		"01100010",
		"01100001",
		"01100000",
		"01100100",
		"01100001",
		"01100011",
		"01101011",
		"01111101",
		"10001110",
		"10011110",
		"10100110",
		"10100101",
		"10001101",
		"01111010",
		"01111101",
		"10000111",
		"10000000",
		"01111010",
		"01110010",
		"01101010",
		"01110101",
		"01110001",
		"01011111",
		"01011101",
		"01100011",
		"01101001",
		"01110011",
		"01101011",
		"01100000",
		"01100011",
		"01110111",
		"01110101",
		"00111011",
		"00010010",
		"00100110",
		"00111010",
		"01001100",
		"01011111",
		"01110011",
		"10000010",
		"10001100",
		"10001110",
		"10011000",
		"10011010",
		"10011110",
		"10100100",
		"10110101",
		"11001010",
		"11010110",
		"11011001",
		"11011001",
		"11010001",
		"10111010",
		"10100110",
		"10100110",
		"10100010",
		"10100010",
		"10001100",
		"01101000",
		"01011110",
		"01010011",
		"01010011",
		"01100010",
		"01111100",
		"10001111",
		"10001111",
		"10010100",
		"10011000",
		"10100000",
		"10100100",
		"10001011",
		"11001010",
		"11000010",
		"11000001",
		"11000011",
		"11000010",
		"10111110",
		"10110011",
		"10011101",
		"01110100",
		"01000000",
		"00100001",
		"00010001",
		"00001110",
		"00010000",
		"00001111",
		"01000100",
		"10101000",
		"10101001",
		"10011111",
		"10011010",
		"10010100",
		"10011000",
		"10100000",
		"10100000",
		"10011110",
		"10100010",
		"10110000",
		"10011010",
		"01111000",
		"10011010",
		"10011111",
		"10001100",
		"10001010",
		"10001101",
		"10001110",
		"10010010",
		"10011100",
		"10011111",
		"10100010",
		"10100110",
		"10100110",
		"10101100",
		"10110001",
		"10111000",
		"10111000",
		"10110000",
		"10101111",
		"10110001",
		"10110011",
		"10110010",
		"10110011",
		"10110111",
		"10111010",
		"10111001",
		"10110101",
		"10111111",
		"10000101",
		"01010100",
		"01011001",
		"01011110",
		"01011110",
		"01100010",
		"01100101",
		"01101011",
		"10001010",
		"11000110",
		"11011001",
		"11011010",
		"10111001",
		"01110010",
		"01100011",
		"01011110",
		"01011100",
		"01010101",
		"01010111",
		"01011001",
		"01011001",
		"01011100",
		"01011110",
		"01100000",
		"01100001",
		"01100000",
		"01011110",
		"01011110",
		"01100001",
		"01101000",
		"01110000",
		"01111011",
		"10000000",
		"01111010",
		"01110101",
		"01111001",
		"01110110",
		"01110101",
		"01110000",
		"01101100",
		"01101011",
		"01101010",
		"01101000",
		"01110011",
		"01100000",
		"01011111",
		"01011101",
		"01100101",
		"10001010",
		"11000100",
		"10111001",
		"01110001",
		"01100011",
		"10000101",
		"01111000",
		"01000000",
		"00010000",
		"00100111",
		"00111101",
		"01010100",
		"01011101",
		"01110001",
		"10000010",
		"10001100",
		"10010001",
		"10011001",
		"10011100",
		"10011101",
		"10101000",
		"10111011",
		"11001110",
		"11010110",
		"11011001",
		"11010111",
		"11001100",
		"10110100",
		"10100010",
		"10100110",
		"10100100",
		"10100001",
		"01111111",
		"01011000",
		"01001101",
		"01011110",
		"10001100",
		"10110100",
		"11010011",
		"10111001",
		"10000100",
		"10001111",
		"10011000",
		"10011101",
		"10100001",
		"01110110",
		"10101000",
		"10100100",
		"10100111",
		"10101011",
		"10101011",
		"10100101",
		"10010101",
		"01111001",
		"01001001",
		"00011011",
		"00001011",
		"00001100",
		"00010011",
		"00010111",
		"00011000",
		"01100110",
		"10101010",
		"10100011",
		"10011000",
		"10001111",
		"10010011",
		"10100000",
		"10011111",
		"10011101",
		"10011101",
		"10100100",
		"10101101",
		"10110010",
		"10010111",
		"10010100",
		"10011001",
		"10010010",
		"10010001",
		"10010001",
		"10010110",
		"10011011",
		"10011110",
		"10100000",
		"10101000",
		"10101100",
		"10101011",
		"10101101",
		"10110010",
		"10111010",
		"10111010",
		"10110001",
		"10110010",
		"10110101",
		"11000000",
		"11001011",
		"11001101",
		"11000101",
		"10111111",
		"10111101",
		"10111000",
		"11000011",
		"10010101",
		"01010010",
		"01011100",
		"01100011",
		"01100010",
		"01100010",
		"01100101",
		"01110000",
		"10001110",
		"11000001",
		"11010111",
		"11011100",
		"11001110",
		"10010011",
		"01100111",
		"01011111",
		"01011011",
		"01010101",
		"01010011",
		"01011000",
		"01011001",
		"01011010",
		"01011101",
		"01011101",
		"01011110",
		"01100000",
		"01100001",
		"01100001",
		"01100010",
		"01100011",
		"01100100",
		"01101100",
		"01110000",
		"01101110",
		"01101110",
		"01110110",
		"01110011",
		"01101110",
		"01101010",
		"01100110",
		"01100100",
		"01100101",
		"01101001",
		"01100000",
		"01011110",
		"01011110",
		"01011101",
		"01101000",
		"10101010",
		"11011100",
		"11100100",
		"10100100",
		"01101001",
		"10010101",
		"10000001",
		"01000010",
		"00010000",
		"00100000",
		"00111101",
		"01010101",
		"01100001",
		"01110010",
		"10001000",
		"10001110",
		"10010001",
		"10010111",
		"10011101",
		"10011111",
		"10101000",
		"10110110",
		"11000101",
		"11010011",
		"11011001",
		"11011000",
		"11001100",
		"10110011",
		"10100001",
		"10100010",
		"10100111",
		"10011101",
		"01100111",
		"01100010",
		"10000100",
		"10111001",
		"11010101",
		"11011101",
		"11000110",
		"10100011",
		"10000011",
		"10010000",
		"10011010",
		"10011100",
		"10100010",
		"01001111",
		"01110101",
		"01110011",
		"01110101",
		"01110111",
		"01111010",
		"01111111",
		"10000101",
		"10001001",
		"10001011",
		"10000011",
		"01101101",
		"01001011",
		"00101011",
		"00011100",
		"00100011",
		"01111101",
		"10100100",
		"10011111",
		"10011010",
		"10001001",
		"10010010",
		"10100000",
		"10011011",
		"10011010",
		"10100000",
		"10100110",
		"10101101",
		"10101011",
		"10001000",
		"10001010",
		"10011000",
		"10011010",
		"10010101",
		"10010011",
		"10010111",
		"10011110",
		"10100011",
		"10101010",
		"10101111",
		"10110000",
		"10101100",
		"10110100",
		"10111000",
		"10111010",
		"10110111",
		"10110000",
		"10110001",
		"10111000",
		"11001011",
		"11011011",
		"11011001",
		"11001011",
		"11000010",
		"10111110",
		"10111011",
		"11000010",
		"10000100",
		"01010011",
		"01100000",
		"01100101",
		"01100011",
		"01100100",
		"01100011",
		"01110100",
		"10010011",
		"10110110",
		"11010011",
		"11011100",
		"11011000",
		"10101110",
		"01110011",
		"01100000",
		"01011100",
		"01010101",
		"01010001",
		"01010111",
		"01011010",
		"01011011",
		"01011011",
		"01011100",
		"01011100",
		"01011101",
		"01011111",
		"01100001",
		"01100010",
		"01100011",
		"01100101",
		"01100111",
		"01101001",
		"01101010",
		"01101100",
		"01101011",
		"01101000",
		"01100110",
		"01100100",
		"01100011",
		"01100011",
		"01100110",
		"01100000",
		"01011101",
		"01011111",
		"01011100",
		"01011110",
		"01111111",
		"10111110",
		"11011001",
		"11011011",
		"10101110",
		"01110011",
		"10001110",
		"01111100",
		"00111001",
		"00010000",
		"00100000",
		"00110110",
		"01001010",
		"01011101",
		"01101101",
		"10000000",
		"10001011",
		"10001100",
		"10010010",
		"10011010",
		"10100011",
		"10101000",
		"10101110",
		"10110001",
		"11000100",
		"11010110",
		"11011010",
		"11010000",
		"10111011",
		"10101001",
		"10011101",
		"10100111",
		"10000000",
		"01110101",
		"10101010",
		"11001010",
		"11011111",
		"11001011",
		"10010001",
		"01101110",
		"01110101",
		"10001010",
		"10010110",
		"10011011",
		"10011111",
		"10100100",
		"01011101",
		"10000110",
		"01111111",
		"01111001",
		"01111011",
		"01111011",
		"10000011",
		"10001001",
		"10010001",
		"10010101",
		"10010101",
		"10010101",
		"10001001",
		"01010000",
		"00010101",
		"00011100",
		"01111110",
		"10011111",
		"10011111",
		"10011001",
		"10001010",
		"10001111",
		"10010010",
		"10001111",
		"10010101",
		"10011101",
		"10100010",
		"10101001",
		"10100010",
		"01111111",
		"10000000",
		"10010110",
		"10100011",
		"10011001",
		"10010100",
		"10010111",
		"10011101",
		"10100100",
		"10101100",
		"10110000",
		"10101100",
		"10110001",
		"10111111",
		"10111111",
		"10111111",
		"10111010",
		"10110001",
		"10110011",
		"10111001",
		"11000111",
		"11010000",
		"11001010",
		"11000000",
		"10111110",
		"10111001",
		"10111001",
		"10111101",
		"01110010",
		"01010100",
		"01100010",
		"01100011",
		"01100001",
		"01100010",
		"01100011",
		"01101100",
		"10001010",
		"10101111",
		"11001100",
		"11011000",
		"11011100",
		"11000110",
		"10000011",
		"01100100",
		"01011110",
		"01010101",
		"01010010",
		"01010111",
		"01011001",
		"01011011",
		"01011001",
		"01011011",
		"01011011",
		"01011011",
		"01011111",
		"01011111",
		"01011111",
		"01100100",
		"01100101",
		"01100110",
		"01101001",
		"01101010",
		"01101000",
		"01100101",
		"01100110",
		"01100101",
		"01100110",
		"01100111",
		"01100101",
		"01011111",
		"01011101",
		"01100000",
		"01011110",
		"01011011",
		"01100101",
		"10011110",
		"11010001",
		"11011001",
		"11001110",
		"10010111",
		"01101101",
		"01110111",
		"01101001",
		"00100101",
		"00010001",
		"00100010",
		"00110100",
		"01000010",
		"01010010",
		"01101001",
		"01111001",
		"10000010",
		"10000100",
		"10001010",
		"10010010",
		"10011100",
		"10100001",
		"10100101",
		"10101000",
		"10110110",
		"11001111",
		"11010111",
		"11010011",
		"11000110",
		"10111001",
		"10100001",
		"10000110",
		"10001110",
		"10111011",
		"11001111",
		"11011011",
		"10110010",
		"01101011",
		"01101000",
		"01111011",
		"10000111",
		"10010000",
		"10010100",
		"10011011",
		"10100010",
		"10100101",
		"01011011",
		"10000101",
		"10010110",
		"10010110",
		"01111100",
		"01110110",
		"10000000",
		"10000111",
		"10001011",
		"10010010",
		"10010001",
		"10001010",
		"01110001",
		"00101011",
		"00001011",
		"00001110",
		"01110110",
		"10100101",
		"10010110",
		"10001111",
		"10001111",
		"10010011",
		"10010010",
		"10001111",
		"10010100",
		"10010110",
		"10011000",
		"10011101",
		"10011001",
		"10000011",
		"01111110",
		"10001101",
		"10100010",
		"10100011",
		"10011010",
		"10011011",
		"10011111",
		"10100011",
		"10101011",
		"10101111",
		"10101110",
		"10111010",
		"11000000",
		"10111111",
		"10111110",
		"10111001",
		"10101110",
		"10101111",
		"10110111",
		"10111100",
		"10111011",
		"10111010",
		"10111011",
		"10111011",
		"10111000",
		"10111000",
		"10111011",
		"10000011",
		"01010000",
		"01011111",
		"01100000",
		"01100000",
		"01100001",
		"01100010",
		"01101001",
		"01111101",
		"10100100",
		"11000011",
		"11010010",
		"11010111",
		"11010001",
		"10011001",
		"01101001",
		"01100011",
		"01011000",
		"01010001",
		"01010010",
		"01010110",
		"01011000",
		"01011010",
		"01011001",
		"01011001",
		"01011010",
		"01011101",
		"01011101",
		"01011110",
		"01100010",
		"01100110",
		"01100110",
		"01101000",
		"01101011",
		"01101001",
		"01101000",
		"01101001",
		"01100111",
		"01100110",
		"01100100",
		"01011111",
		"01011110",
		"01100011",
		"01100000",
		"01011101",
		"01011111",
		"01111110",
		"10111111",
		"11010110",
		"11001110",
		"10101111",
		"01110100",
		"01100101",
		"01100111",
		"01010010",
		"00010010",
		"00010100",
		"00100101",
		"00111000",
		"01000100",
		"01001001",
		"01011011",
		"01110001",
		"01110110",
		"01111011",
		"10000000",
		"10000101",
		"10001111",
		"10011011",
		"10100011",
		"10100001",
		"10110111",
		"11001110",
		"11001111",
		"11001110",
		"11000100",
		"10110100",
		"10001011",
		"10010010",
		"10111100",
		"11010000",
		"11011000",
		"10011111",
		"01010011",
		"01100001",
		"01110100",
		"10000000",
		"10001000",
		"10001011",
		"10010100",
		"10011110",
		"10100001",
		"10100100",
		"01010010",
		"01101111",
		"10001000",
		"10101010",
		"10100111",
		"10001010",
		"01111000",
		"01111101",
		"10000010",
		"10001001",
		"10001010",
		"01110111",
		"00111111",
		"00001110",
		"00001001",
		"00001110",
		"01010011",
		"10011001",
		"10011000",
		"10001011",
		"10010101",
		"10010101",
		"10001101",
		"10001010",
		"10001110",
		"10001101",
		"10001010",
		"10001100",
		"10001100",
		"10001100",
		"10000001",
		"10001000",
		"10010111",
		"10100011",
		"10011110",
		"10011011",
		"10100000",
		"10100100",
		"10101010",
		"10101100",
		"10101111",
		"10110111",
		"10111011",
		"10111011",
		"10111011",
		"10110111",
		"10101110",
		"10101110",
		"10110010",
		"10110011",
		"10111000",
		"10111010",
		"10111011",
		"10111010",
		"10111001",
		"10111001",
		"10111011",
		"10100010",
		"01010110",
		"01011011",
		"01011111",
		"01100000",
		"01100000",
		"01100000",
		"01100110",
		"01110101",
		"10001101",
		"10100001",
		"10101011",
		"10110010",
		"10110001",
		"10010010",
		"01101111",
		"01100111",
		"01100000",
		"01010010",
		"01001100",
		"01001011",
		"01010101",
		"01011001",
		"01010111",
		"01010110",
		"01010011",
		"01010110",
		"01011011",
		"01011110",
		"01100000",
		"01100100",
		"01100101",
		"01100101",
		"01100111",
		"01101000",
		"01101000",
		"01100101",
		"01100010",
		"01011110",
		"01011110",
		"01100001",
		"01100100",
		"01100011",
		"01100001",
		"01101001",
		"10000101",
		"10110000",
		"11001001",
		"10111010",
		"10010100",
		"01110111",
		"01100100",
		"01100000",
		"01100011",
		"00110001",
		"00001011",
		"00010100",
		"00100010",
		"00111000",
		"01000001",
		"01000110",
		"01010001",
		"01100000",
		"01101011",
		"01110010",
		"01111010",
		"10000010",
		"10000011",
		"10010001",
		"10010111",
		"10010110",
		"10101011",
		"11000000",
		"11000110",
		"10111111",
		"10101111",
		"10010001",
		"10001111",
		"10111010",
		"11001011",
		"11010101",
		"10111001",
		"01000100",
		"01001001",
		"01011001",
		"01100110",
		"01110100",
		"10000000",
		"10001001",
		"10010100",
		"10011010",
		"10011111",
		"10100010",
		"01010000",
		"01011011",
		"01011100",
		"01110101",
		"10010111",
		"10011101",
		"01110110",
		"01101100",
		"01110011",
		"01110001",
		"01011110",
		"00110011",
		"00001111",
		"00001000",
		"00001001",
		"00011010",
		"01001011",
		"10000001",
		"10010010",
		"10000110",
		"10001010",
		"10001010",
		"10001001",
		"10000111",
		"10000010",
		"10000001",
		"10000011",
		"10000001",
		"01111101",
		"10001010",
		"10001011",
		"10001000",
		"10010010",
		"10011010",
		"10011010",
		"10011001",
		"10011010",
		"10011111",
		"10100011",
		"10101010",
		"10101101",
		"10101111",
		"10110000",
		"10110001",
		"10110101",
		"10110110",
		"10110010",
		"10110001",
		"10110011",
		"10110101",
		"10111001",
		"10111010",
		"10111010",
		"10111011",
		"10111001",
		"10111001",
		"10111001",
		"10110001",
		"01011001",
		"01010101",
		"01011110",
		"01011110",
		"01011111",
		"01100000",
		"01100011",
		"01101100",
		"01110111",
		"01111110",
		"01111001",
		"10000010",
		"10001001",
		"10000001",
		"01110011",
		"01101011",
		"01100110",
		"01011100",
		"01010101",
		"01001010",
		"01000011",
		"01010000",
		"01010111",
		"01011000",
		"01011111",
		"01100101",
		"01010100",
		"01011000",
		"01100000",
		"01100000",
		"01100001",
		"01100001",
		"01100001",
		"01100001",
		"01100001",
		"01100001",
		"01100011",
		"01100000",
		"01100001",
		"01100001",
		"01100100",
		"01100010",
		"01101010",
		"10010111",
		"10111110",
		"11001110",
		"10111110",
		"10010000",
		"01110001",
		"01100110",
		"01100000",
		"01011101",
		"01010111",
		"00010101",
		"00001010",
		"00010001",
		"00011010",
		"00101011",
		"00111000",
		"00111110",
		"01000100",
		"01001001",
		"01001100",
		"01010110",
		"01100011",
		"01100101",
		"01100101",
		"01101100",
		"01110010",
		"01111001",
		"01110010",
		"01111111",
		"01111110",
		"01101110",
		"01111010",
		"10001100",
		"10101100",
		"11001100",
		"11010011",
		"11010101",
		"10111111",
		"10100011",
		"10100110",
		"10011010",
		"01111011",
		"01100111",
		"01101110",
		"10000000",
		"10001101",
		"10010011",
		"10011101",
		"10100000",
		"00110110",
		"01010001",
		"01010010",
		"01010000",
		"01001110",
		"01001110",
		"01001010",
		"01000100",
		"01000010",
		"00111000",
		"00011100",
		"00001001",
		"00001000",
		"00001000",
		"00000111",
		"00010000",
		"01011011",
		"10001101",
		"10010101",
		"10000101",
		"10000101",
		"10000110",
		"10000000",
		"01111011",
		"01110001",
		"01101011",
		"01100000",
		"01010000",
		"01001110",
		"10001010",
		"10010011",
		"10001100",
		"10001111",
		"10010011",
		"10010101",
		"10010110",
		"10010111",
		"10011101",
		"10100100",
		"10101010",
		"10101110",
		"10101100",
		"10101111",
		"10110000",
		"10110011",
		"10110110",
		"10110110",
		"10110101",
		"10110110",
		"10110111",
		"10111011",
		"10111010",
		"10111010",
		"10111011",
		"10111010",
		"10111011",
		"10111001",
		"10110010",
		"01010110",
		"01010010",
		"01011010",
		"01011110",
		"01011111",
		"01011110",
		"01011111",
		"01100101",
		"01101001",
		"01110001",
		"01110011",
		"01110110",
		"01111010",
		"01111001",
		"01110110",
		"01101111",
		"01101000",
		"01100100",
		"01101010",
		"01110101",
		"10000000",
		"10001000",
		"10010101",
		"10100110",
		"10110111",
		"10101100",
		"10001110",
		"01011111",
		"01010000",
		"01010111",
		"01011010",
		"01011101",
		"01011101",
		"01011101",
		"01100001",
		"01100001",
		"01100011",
		"01100100",
		"01100011",
		"01100010",
		"01100100",
		"01101011",
		"10001001",
		"10110011",
		"11000100",
		"11000011",
		"10100101",
		"01111011",
		"01101000",
		"01100010",
		"01011101",
		"01011110",
		"00111010",
		"00000001",
		"00001001",
		"00010000",
		"00010110",
		"00011111",
		"00101000",
		"00101101",
		"00110000",
		"00110000",
		"00110010",
		"00110110",
		"00101100",
		"00100001",
		"00110000",
		"01100110",
		"10001001",
		"10010011",
		"01011110",
		"01001000",
		"01101110",
		"10011100",
		"10110111",
		"10100101",
		"11000000",
		"11001110",
		"11010011",
		"11010010",
		"11010001",
		"11010000",
		"11001010",
		"11000100",
		"11001001",
		"11000100",
		"10100010",
		"01111111",
		"10000011",
		"10001100",
		"10011000",
		"10011101",
		"00100011",
		"00101101",
		"00110001",
		"00101001",
		"00011111",
		"00011100",
		"00011111",
		"00011000",
		"00010001",
		"00001100",
		"00000110",
		"00000011",
		"00000010",
		"00001010",
		"00011010",
		"00101010",
		"01011010",
		"01100011",
		"01011001",
		"01001100",
		"01100011",
		"10000100",
		"01111000",
		"01100000",
		"01001100",
		"00110110",
		"00101100",
		"00100001",
		"00110010",
		"10001111",
		"10010011",
		"10010000",
		"10010001",
		"10011000",
		"10010110",
		"10011001",
		"10010111",
		"10011000",
		"10100000",
		"10100101",
		"10101001",
		"10101010",
		"10101100",
		"10101111",
		"10110011",
		"10111001",
		"10111011",
		"11000000",
		"11000011",
		"10111101",
		"10111011",
		"10111000",
		"10111001",
		"10111010",
		"10111001",
		"10111010",
		"10110111",
		"10101011",
		"01001101",
		"01010000",
		"01011000",
		"01011100",
		"01011100",
		"01011101",
		"01011110",
		"01011111",
		"01100001",
		"01100110",
		"01100110",
		"01101010",
		"01101101",
		"01110011",
		"01110010",
		"01101110",
		"01101100",
		"01101110",
		"01110100",
		"01111100",
		"01111111",
		"01111100",
		"10001010",
		"10110111",
		"11000111",
		"11000111",
		"11000111",
		"10100100",
		"01001000",
		"01010001",
		"01011000",
		"01011110",
		"01011111",
		"01100000",
		"01100010",
		"01100001",
		"01100000",
		"01100001",
		"01100001",
		"01100100",
		"01101001",
		"01111111",
		"10101010",
		"10111111",
		"10111000",
		"10011010",
		"01111010",
		"01101001",
		"01100011",
		"01011111",
		"01011101",
		"01011101",
		"01000110",
		"01011111",
		"01000000",
		"00001001",
		"00001111",
		"00010011",
		"00010011",
		"00010111",
		"00011100",
		"00100001",
		"00011101",
		"00010111",
		"00001001",
		"00110101",
		"10011000",
		"10111101",
		"11000001",
		"10101111",
		"10100001",
		"10100010",
		"10100111",
		"10101110",
		"10111001",
		"10111000",
		"11001110",
		"11001100",
		"11010001",
		"11010001",
		"11001101",
		"11001011",
		"11001010",
		"11000101",
		"11001111",
		"11010111",
		"11011001",
		"11000001",
		"01111110",
		"10000000",
		"10010000",
		"10010100",
		"00010010",
		"00001101",
		"00010011",
		"00001111",
		"00001101",
		"00001100",
		"00001011",
		"00001011",
		"00001000",
		"00000010",
		"00000101",
		"00100100",
		"01010001",
		"01100110",
		"01011001",
		"01000011",
		"00110001",
		"00100010",
		"00011011",
		"00110110",
		"01100101",
		"01101001",
		"01011001",
		"01000110",
		"00110111",
		"00110100",
		"00110100",
		"00101000",
		"01001010",
		"10011011",
		"10010011",
		"10010000",
		"10010010",
		"10011000",
		"10010111",
		"10011000",
		"10011001",
		"10011010",
		"10100000",
		"10100011",
		"10100100",
		"10100101",
		"10101010",
		"10101110",
		"10110000",
		"10110111",
		"10111110",
		"11000100",
		"11000001",
		"10111100",
		"10111010",
		"10111001",
		"10111011",
		"10111011",
		"10111001",
		"10111001",
		"10110110",
		"10100000",
		"01000111",
		"01001100",
		"01010101",
		"01011001",
		"01011011",
		"01011011",
		"01011100",
		"01011111",
		"01100001",
		"01100010",
		"01100010",
		"01100100",
		"01101001",
		"01101100",
		"01101101",
		"01101110",
		"01101100",
		"01101001",
		"01100011",
		"01010101",
		"01010100",
		"01011001",
		"01101000",
		"10001011",
		"10111101",
		"11001000",
		"10111001",
		"11001100",
		"01101001",
		"01001011",
		"01011001",
		"01011110",
		"01100011",
		"01100010",
		"01100011",
		"01100010",
		"01100010",
		"01100101",
		"01100111",
		"01101010",
		"01110111",
		"10000110",
		"10010111",
		"10100110",
		"10011111",
		"10000100",
		"01110001",
		"01100011",
		"01100000",
		"01011101",
		"01011110",
		"01100111",
		"10011001",
		"10101000",
		"00100111",
		"00001001",
		"00001111",
		"00001111",
		"00001101",
		"00001111",
		"00010000",
		"00001111",
		"00001110",
		"00000111",
		"00100101",
		"10011101",
		"10111000",
		"10111001",
		"10111000",
		"10110100",
		"10111100",
		"10111101",
		"10101101",
		"10110100",
		"10101001",
		"10110010",
		"11001110",
		"11000111",
		"11001100",
		"11001100",
		"11000110",
		"11000011",
		"11000011",
		"11001111",
		"11010101",
		"11010101",
		"11010100",
		"11011010",
		"10101100",
		"01110001",
		"10000110",
		"10001110",
		"01001101",
		"01010001",
		"00111101",
		"00100101",
		"00010001",
		"00000110",
		"00000100",
		"00000001",
		"00001010",
		"00111000",
		"01110011",
		"10000010",
		"01100001",
		"01000000",
		"00110001",
		"00110000",
		"00101011",
		"00101011",
		"01000010",
		"01100100",
		"01100101",
		"01010101",
		"01000011",
		"00110101",
		"00110010",
		"00110000",
		"00101110",
		"00100111",
		"01011111",
		"10100000",
		"10011000",
		"10010001",
		"10010001",
		"10010111",
		"10010101",
		"10010110",
		"10011000",
		"10011100",
		"10100000",
		"10100011",
		"10100111",
		"10100110",
		"10101010",
		"10101101",
		"10110011",
		"10110110",
		"10111011",
		"11000001",
		"10111101",
		"10111100",
		"10111011",
		"10111100",
		"10111110",
		"10111100",
		"10111011",
		"10111010",
		"10110111",
		"10010010",
		"01000100",
		"01001101",
		"01010011",
		"01010111",
		"01010111",
		"01010111",
		"01011001",
		"01011101",
		"01100000",
		"01100001",
		"01100001",
		"01100011",
		"01100111",
		"01101111",
		"01110001",
		"01101101",
		"01101011",
		"01101011",
		"01101010",
		"01101011",
		"01011100",
		"01010000",
		"01101001",
		"01110011",
		"10100010",
		"11001000",
		"11000001",
		"11000100",
		"10100111",
		"01001100",
		"01010011",
		"01011001",
		"01011110",
		"01100000",
		"01100010",
		"01100000",
		"01100011",
		"01100110",
		"01101000",
		"01101101",
		"01111101",
		"10000110",
		"10000100",
		"10000011",
		"01111110",
		"01110011",
		"01101010",
		"01100010",
		"01100010",
		"01100000",
		"01011111",
		"01100011",
		"10100100",
		"10101111",
		"00011110",
		"00000110",
		"00001100",
		"00001101",
		"00001101",
		"00001100",
		"00001011",
		"00001101",
		"00001100",
		"00001010",
		"01101001",
		"10110000",
		"10110011",
		"10110101",
		"10110111",
		"10111111",
		"11000011",
		"11001000",
		"11001001",
		"11000101",
		"10111100",
		"10111110",
		"11000111",
		"11001001",
		"11001101",
		"11001111",
		"11010000",
		"11010001",
		"11010000",
		"11010011",
		"11010100",
		"11010101",
		"11010101",
		"11010111",
		"11000010",
		"01101101",
		"01111110",
		"10001000",
		"01101111",
		"10010110",
		"10001101",
		"10000110",
		"01110111",
		"01011101",
		"00110111",
		"00101101",
		"01110110",
		"10010011",
		"01111000",
		"01001111",
		"00110110",
		"00101110",
		"00101110",
		"00101101",
		"00101001",
		"01000010",
		"01101000",
		"01100011",
		"01010011",
		"01000001",
		"00110100",
		"00101111",
		"00110001",
		"00101111",
		"00101100",
		"00100110",
		"01110000",
		"10011110",
		"10011011",
		"10010110",
		"10010000",
		"10010101",
		"10010101",
		"10010110",
		"10011000",
		"10011010",
		"10100000",
		"10100010",
		"10100100",
		"10100100",
		"10101000",
		"10101111",
		"10110101",
		"10111001",
		"10111011",
		"10111100",
		"10111101",
		"10111100",
		"10111100",
		"10111100",
		"10111111",
		"10111111",
		"10111110",
		"10111010",
		"10110110",
		"01111111",
		"01000011",
		"01001101",
		"01010010",
		"01010010",
		"01010011",
		"01010110",
		"01011001",
		"01011100",
		"01011101",
		"01011110",
		"01011110",
		"01100000",
		"01100010",
		"01100111",
		"01101001",
		"01101011",
		"01101101",
		"01101100",
		"01101100",
		"01101000",
		"01100100",
		"01010011",
		"01110111",
		"01111110",
		"10001001",
		"10111010",
		"11001010",
		"10111011",
		"11010010",
		"01110010",
		"01000100",
		"01010010",
		"01010111",
		"01011000",
		"01011100",
		"01011101",
		"01011110",
		"01100001",
		"01100011",
		"01100100",
		"01101001",
		"01101011",
		"01101001",
		"01100110",
		"01100010",
		"01100001",
		"01100010",
		"01100110",
		"01101010",
		"01100110",
		"01000111",
		"00101000",
		"10000111",
		"10011010",
		"01001011",
		"00001000",
		"00000110",
		"00001010",
		"00001001",
		"00001010",
		"00001100",
		"00001101",
		"00001001",
		"00010101",
		"10001000",
		"10101101",
		"10101111",
		"10110010",
		"10110110",
		"10111110",
		"11000110",
		"11001000",
		"11001001",
		"11001001",
		"11000111",
		"11000111",
		"11001001",
		"11001101",
		"11010000",
		"11010010",
		"11010101",
		"11010110",
		"11010110",
		"11010101",
		"11010100",
		"11010100",
		"11010101",
		"11011000",
		"10111101",
		"01100001",
		"01110101",
		"01111110",
		"01110010",
		"10011100",
		"10010100",
		"10001111",
		"10000111",
		"01101110",
		"01110000",
		"10001010",
		"01111110",
		"01100011",
		"01010001",
		"00111111",
		"00110101",
		"00110100",
		"00110010",
		"00110000",
		"00110110",
		"01010101",
		"01011011",
		"01001101",
		"00111101",
		"00110010",
		"00110001",
		"00110000",
		"00110011",
		"00110000",
		"00101010",
		"00101101",
		"10000110",
		"10011001",
		"10011110",
		"10100000",
		"10011001",
		"10010010",
		"10010011",
		"10010100",
		"10010111",
		"10011000",
		"10011011",
		"10100010",
		"10100011",
		"10100001",
		"10101011",
		"10110010",
		"10111000",
		"10111010",
		"10111011",
		"10111101",
		"10111111",
		"10111011",
		"10111011",
		"10111100",
		"10111110",
		"11000000",
		"10111110",
		"10110111",
		"10110101",
		"01101110",
		"00111111",
		"01001000",
		"01001110",
		"01010001",
		"01010011",
		"01010101",
		"01011000",
		"01011011",
		"01011100",
		"01011110",
		"01011111",
		"01100000",
		"01100100",
		"01101000",
		"01101010",
		"01101101",
		"01101110",
		"01101100",
		"01100111",
		"01100010",
		"01011101",
		"01001111",
		"01101101",
		"10000011",
		"01111011",
		"10100110",
		"11000111",
		"10111100",
		"11000001",
		"10110011",
		"01000111",
		"01001000",
		"01001111",
		"01010110",
		"01011001",
		"01011010",
		"01011100",
		"01011110",
		"01011110",
		"01011100",
		"01011100",
		"01011100",
		"01011011",
		"01011110",
		"01100001",
		"01100011",
		"01100111",
		"01101101",
		"01101010",
		"01000110",
		"00001100",
		"00000111",
		"00100101",
		"01000100",
		"01100110",
		"01001001",
		"00001110",
		"00000100",
		"00000100",
		"00000101",
		"00001001",
		"00001010",
		"00001000",
		"00011000",
		"10001100",
		"10101000",
		"10101001",
		"10101101",
		"10110010",
		"10111010",
		"11000010",
		"11000110",
		"11000110",
		"11000110",
		"11000110",
		"11001000",
		"11001010",
		"11001101",
		"11010000",
		"11010011",
		"11010101",
		"11011000",
		"11011001",
		"11011001",
		"11010110",
		"11010101",
		"11010101",
		"11011011",
		"10101111",
		"01010010",
		"01101001",
		"01110110",
		"01110101",
		"10011101",
		"10010110",
		"10010101",
		"01111011",
		"01101101",
		"10000110",
		"01111100",
		"01011111",
		"01001111",
		"01000011",
		"00110111",
		"00110010",
		"00110001",
		"00110011",
		"00110110",
		"01000111",
		"01010011",
		"01000110",
		"00111011",
		"00110101",
		"00110101",
		"00110100",
		"00110010",
		"00110011",
		"00110001",
		"00101010",
		"00111111",
		"10011001",
		"10011111",
		"10011101",
		"10100110",
		"10100001",
		"10011000",
		"10010011",
		"10010100",
		"10010100",
		"10010101",
		"10011000",
		"10011101",
		"10011111",
		"10100011",
		"10101100",
		"10110001",
		"10110110",
		"10111011",
		"10111100",
		"10111101",
		"10111111",
		"10111011",
		"10111011",
		"10111011",
		"10111110",
		"10111110",
		"10111100",
		"10110101",
		"10110011",
		"01100011",
		"00111100",
		"01000100",
		"01001010",
		"01001100",
		"01001111",
		"01010011",
		"01011000",
		"01011010",
		"01011101",
		"01011111",
		"01100010",
		"01100010",
		"01100101",
		"01100111",
		"01101001",
		"01101001",
		"01100101",
		"01100000",
		"01100100",
		"01101010",
		"01100111",
		"01100110",
		"01110000",
		"10001010",
		"01111011",
		"10010001",
		"10110110",
		"11001010",
		"10101101",
		"11010010",
		"01101111",
		"00111110",
		"01001010",
		"01010001",
		"01010010",
		"01010110",
		"01011011",
		"01100000",
		"01100101",
		"01101000",
		"01100100",
		"01100100",
		"01100111",
		"01100100",
		"01011100",
		"01011000",
		"01011001",
		"01011010",
		"00110110",
		"00001111",
		"00011101",
		"01000110",
		"01101110",
		"10000101",
		"10000000",
		"10000001",
		"01100010",
		"01000011",
		"00101111",
		"00011000",
		"00001000",
		"00000111",
		"00000111",
		"00011001",
		"10001010",
		"10100100",
		"10100100",
		"10100111",
		"10101100",
		"10110101",
		"10111011",
		"10111111",
		"10111101",
		"11000000",
		"11000010",
		"11000011",
		"11000110",
		"11001100",
		"11001111",
		"11010001",
		"11010100",
		"11010110",
		"11010110",
		"11010110",
		"11010110",
		"11010101",
		"11010100",
		"11011100",
		"10010011",
		"00111111",
		"01100000",
		"01110010",
		"01110100",
		"10011010",
		"10010010",
		"01110101",
		"01101011",
		"10000011",
		"01111100",
		"01101000",
		"01010110",
		"01001001",
		"00111100",
		"00111000",
		"00110101",
		"00110100",
		"00110111",
		"00111110",
		"01000111",
		"01000011",
		"00111001",
		"00110100",
		"00110110",
		"00110100",
		"00110101",
		"00110011",
		"00110000",
		"00110000",
		"00100101",
		"01010100",
		"10011111",
		"10100111",
		"10100011",
		"10100110",
		"10100000",
		"10011111",
		"10011011",
		"10011000",
		"10010110",
		"10010100",
		"10011000",
		"10011010",
		"10011101",
		"10100101",
		"10101100",
		"10101111",
		"10110101",
		"10111010",
		"10111010",
		"10111101",
		"10111011",
		"10111010",
		"10111100",
		"10111101",
		"10111100",
		"10111001",
		"10111011",
		"10110110",
		"10110011",
		"01011010",
		"00110111",
		"01000000",
		"01000100",
		"01000111",
		"01001100",
		"01001101",
		"01010100",
		"01011001",
		"01100010",
		"01011011",
		"01011100",
		"01011101",
		"01011111",
		"01011111",
		"01011010",
		"01010001",
		"01010000",
		"01101001",
		"01111010",
		"10000011",
		"10010000",
		"10011011",
		"10010101",
		"10000110",
		"10001111",
		"10001000",
		"10100111",
		"11001110",
		"10110001",
		"11000100",
		"10101101",
		"01000101",
		"01000110",
		"01000100",
		"01001011",
		"01011100",
		"01101011",
		"01111011",
		"01111101",
		"01110101",
		"01111110",
		"10001101",
		"10011101",
		"10100101",
		"10011010",
		"10000100",
		"01101001",
		"00100111",
		"00000111",
		"00100101",
		"01101000",
		"10010111",
		"10011111",
		"10100001",
		"10100010",
		"10100001",
		"10100000",
		"10010111",
		"10001000",
		"01110010",
		"01001000",
		"00010110",
		"00000101",
		"00001110",
		"01111001",
		"10011110",
		"10100000",
		"10100011",
		"10100100",
		"10101110",
		"10110110",
		"10111010",
		"10111010",
		"10111101",
		"10111111",
		"11000000",
		"11000011",
		"11001000",
		"11001011",
		"11001110",
		"11010011",
		"11010100",
		"11010101",
		"11010110",
		"11010110",
		"11010110",
		"11010110",
		"11011011",
		"01100110",
		"00101110",
		"01011010",
		"01101001",
		"01110111",
		"10001100",
		"01101010",
		"01101110",
		"10000011",
		"01111100",
		"01100110",
		"01010010",
		"01000010",
		"00111010",
		"00110111",
		"00110111",
		"00111000",
		"00111000",
		"00111000",
		"00111010",
		"00111110",
		"00111001",
		"00110110",
		"00110110",
		"00110011",
		"00110010",
		"00110001",
		"00110011",
		"00110000",
		"00101100",
		"00100010",
		"01101000",
		"10011101",
		"10101000",
		"10101001",
		"10100110",
		"10100001",
		"10011111",
		"10100000",
		"10100000",
		"10011110",
		"10011100",
		"10011100",
		"10011101",
		"10011111",
		"10100111",
		"10101100",
		"10110000",
		"10110101",
		"10111000",
		"10111010",
		"10111100",
		"10111011",
		"10111100",
		"10111110",
		"10111110",
		"10111011",
		"10111011",
		"10111100",
		"10110100",
		"10110001",
		"01001001",
		"00110100",
		"00111101",
		"01000001",
		"01000100",
		"01000100",
		"01000110",
		"01000111",
		"01001011",
		"01001101",
		"01001011",
		"01001001",
		"01001010",
		"01001001",
		"01000000",
		"00111010",
		"01001010",
		"01101100",
		"01111110",
		"10001000",
		"10010010",
		"10011110",
		"10100011",
		"10101111",
		"10001010",
		"10001011",
		"10001001",
		"10011011",
		"11000110",
		"11000000",
		"10110010",
		"11010001",
		"01111111",
		"01001000",
		"01001100",
		"01011010",
		"01100111",
		"01111100",
		"01110011",
		"01100000",
		"01100101",
		"01111001",
		"10010110",
		"10011011",
		"10011010",
		"10011111",
		"10101000",
		"10101100",
		"10001110",
		"01010011",
		"01000001",
		"01110111",
		"10010101",
		"10011101",
		"10011111",
		"10100001",
		"10100101",
		"10100100",
		"10100000",
		"10011011",
		"10010100",
		"10000000",
		"01011000",
		"00011111",
		"00000110",
		"01101000",
		"10011000",
		"10011001",
		"10011011",
		"10100000",
		"10100110",
		"10101100",
		"10110010",
		"10110101",
		"10110111",
		"10111001",
		"10111011",
		"10111110",
		"11000001",
		"11000100",
		"11001001",
		"11010000",
		"11010011",
		"11010100",
		"11010101",
		"11010101",
		"11010100",
		"11011000",
		"11000101",
		"00101011",
		"00010001",
		"00101000",
		"01000000",
		"01011111",
		"01110100",
		"01110010",
		"01110111",
		"01110110",
		"01100100",
		"01001011",
		"00111011",
		"00110101",
		"00101111",
		"00101111",
		"00110100",
		"00110100",
		"00110011",
		"00110101",
		"00111001",
		"00111010",
		"00111000",
		"00110111",
		"00110100",
		"00110101",
		"00110101",
		"00110011",
		"00110010",
		"00110010",
		"00101101",
		"00101000",
		"10000100",
		"10011100",
		"10100110",
		"10100111",
		"10100101",
		"10100001",
		"10011111",
		"10100000",
		"10100000",
		"10011100",
		"10011100",
		"10011110",
		"10011111",
		"10100100",
		"10101010",
		"10101101",
		"10110011",
		"10110111",
		"10110111",
		"10111010",
		"10111011",
		"10111100",
		"10111100",
		"10111010",
		"10111100",
		"10111100",
		"10111101",
		"10111011",
		"10110101",
		"10100100",
		"00101111",
		"00100110",
		"00101110",
		"00110000",
		"00101111",
		"00101101",
		"00110000",
		"00101101",
		"00101101",
		"00101111",
		"00110010",
		"00111001",
		"00111111",
		"00101111",
		"00110110",
		"01010001",
		"01110111",
		"10001111",
		"10010001",
		"10010010",
		"10010010",
		"10011101",
		"10101000",
		"10101111",
		"10001110",
		"10000110",
		"10000100",
		"10000101",
		"10110110",
		"11000100",
		"10110000",
		"11001011",
		"10111001",
		"01010100",
		"01010010",
		"01100000",
		"01110001",
		"01110010",
		"01011111",
		"01011010",
		"01101000",
		"10000010",
		"10001100",
		"10010101",
		"10011110",
		"10100010",
		"10100001",
		"10100100",
		"10101011",
		"10101101",
		"10011100",
		"10000011",
		"10000101",
		"10011010",
		"10100001",
		"10100110",
		"10100111",
		"10100100",
		"10100010",
		"10100001",
		"10011110",
		"10010100",
		"10000010",
		"01010000",
		"00001110",
		"01000011",
		"10001110",
		"10010100",
		"10010111",
		"10011100",
		"10100000",
		"10100100",
		"10101001",
		"10101101",
		"10110001",
		"10110100",
		"10110111",
		"10111010",
		"10111100",
		"10111110",
		"11000011",
		"11001010",
		"11001111",
		"11010000",
		"11010001",
		"11010000",
		"11010000",
		"11010100",
		"10000010",
		"00001100",
		"00111001",
		"01110001",
		"01100111",
		"01010100",
		"01111001",
		"01111000",
		"01110100",
		"01100001",
		"01001101",
		"01000000",
		"00110100",
		"00110011",
		"00110001",
		"00101111",
		"00110010",
		"00101101",
		"00110011",
		"00110111",
		"00111001",
		"00111001",
		"00111000",
		"00110101",
		"00110100",
		"00110100",
		"00110011",
		"00110011",
		"00110001",
		"00110010",
		"00101110",
		"01000011",
		"10010111",
		"10100011",
		"10101010",
		"10101000",
		"10100011",
		"10011111",
		"10011110",
		"10100000",
		"10011110",
		"10011101",
		"10011111",
		"10100001",
		"10100100",
		"10101011",
		"10101110",
		"10110000",
		"10110110",
		"10111000",
		"10111001",
		"10111100",
		"10111011",
		"10111011",
		"10111010",
		"10111011",
		"10111110",
		"10111110",
		"10111110",
		"10111001",
		"10111010",
		"10001100",
		"00011010",
		"00011011",
		"00011110",
		"00100001",
		"00100001",
		"00100011",
		"00101101",
		"00111100",
		"01001100",
		"01010111",
		"01011101",
		"01100100",
		"01100000",
		"01010110",
		"01110011",
		"10001101",
		"10001100",
		"10001110",
		"10011110",
		"10100110",
		"10011101",
		"10011010",
		"10100111",
		"10101110",
		"10010111",
		"10000111",
		"10010000",
		"10000001",
		"10100001",
		"10111011",
		"10111011",
		"11000010",
		"11010010",
		"01111111",
		"01000101",
		"01011100",
		"01101000",
		"01011111",
		"01011000",
		"01100001",
		"01110110",
		"01111011",
		"10000101",
		"10010100",
		"10011001",
		"10100000",
		"10100110",
		"10101011",
		"10101111",
		"10110000",
		"10110010",
		"10101110",
		"10011011",
		"10010101",
		"10011110",
		"10100110",
		"10101011",
		"10101101",
		"10101110",
		"10110010",
		"10101111",
		"10011110",
		"10010011",
		"01110100",
		"00101001",
		"00011001",
		"01101010",
		"10000111",
		"10010010",
		"10011000",
		"10011000",
		"10011011",
		"10100001",
		"10100101",
		"10100110",
		"10101100",
		"10101110",
		"10110010",
		"10110011",
		"10111000",
		"10111101",
		"11000011",
		"11000110",
		"11000110",
		"11000101",
		"11000011",
		"10111110",
		"10110001",
		"01110101",
		"10011011",
		"10111000",
		"10010011",
		"01010011",
		"01011011",
		"01111110",
		"01111010",
		"01100100",
		"01010000",
		"01000110",
		"00111110",
		"00110110",
		"00110011",
		"00110001",
		"00110000",
		"00110010",
		"00110001",
		"00110011",
		"00110101",
		"00111000",
		"00111000",
		"00110101",
		"00110011",
		"00110010",
		"00110011",
		"00110001",
		"00110000",
		"00110010",
		"00110000",
		"00101011",
		"01100100",
		"10011100",
		"10101000",
		"10101001",
		"10100111",
		"10100100",
		"10011111",
		"10011111",
		"10100001",
		"10100000",
		"10011111",
		"10100001",
		"10100100",
		"10101000",
		"10101101",
		"10110000",
		"10110011",
		"10110111",
		"10111011",
		"10111010",
		"10111110",
		"10111101",
		"10111011",
		"10111010",
		"10111101",
		"10111111",
		"10111111",
		"10111110",
		"10110111",
		"10110111",
		"01110001",
		"00110001",
		"00110111",
		"00110011",
		"00110010",
		"00111111",
		"01011010",
		"01101101",
		"01111000",
		"10000000",
		"10000100",
		"10000110",
		"10000100",
		"01110101",
		"01011110",
		"01010111",
		"01110001",
		"10010001",
		"10001110",
		"01110100",
		"01101011",
		"10000101",
		"10101010",
		"10110101",
		"10111110",
		"10100001",
		"01111010",
		"10001110",
		"01111110",
		"10001110",
		"10101111",
		"11000001",
		"10111011",
		"11001101",
		"10111111",
		"01011100",
		"01011110",
		"10011101",
		"01110010",
		"01001110",
		"01100001",
		"01110100",
		"01111110",
		"10000101",
		"10001010",
		"10010101",
		"10100010",
		"10101000",
		"10110000",
		"10110111",
		"10111000",
		"10110011",
		"10101100",
		"10101101",
		"10100110",
		"10011111",
		"10100101",
		"10101010",
		"10111000",
		"11000101",
		"11001101",
		"11001100",
		"10110111",
		"10100000",
		"10001100",
		"01010001",
		"00010001",
		"00110100",
		"01100111",
		"01110101",
		"10000100",
		"10001110",
		"10010010",
		"10010100",
		"10010111",
		"10011010",
		"10011110",
		"10011111",
		"10100001",
		"10100001",
		"10100110",
		"10101010",
		"10101110",
		"10110000",
		"10101110",
		"10101000",
		"10100111",
		"10101000",
		"10110011",
		"10101110",
		"10001001",
		"01011111",
		"01001111",
		"01000101",
		"01011100",
		"01111010",
		"01101010",
		"01011000",
		"01001100",
		"01000101",
		"00111100",
		"00110101",
		"00110101",
		"00110011",
		"00110011",
		"00110101",
		"00110100",
		"00110101",
		"00110110",
		"00110110",
		"00110110",
		"00110111",
		"00110110",
		"00110011",
		"00110011",
		"00110010",
		"00110001",
		"00110010",
		"00110000",
		"00101011",
		"01111100",
		"10011110",
		"10101001",
		"10101001",
		"10100100",
		"10100010",
		"10011111",
		"10100000",
		"10100010",
		"10100001",
		"10100010",
		"10100100",
		"10100111",
		"10101010",
		"10101101",
		"10110001",
		"10110110",
		"10111010",
		"10111100",
		"10111010",
		"11000000",
		"10111101",
		"10111011",
		"10111100",
		"10111111",
		"11000001",
		"11000000",
		"10111111",
		"10110101",
		"10101100",
		"01010010",
		"00110111",
		"00111010",
		"01000000",
		"01100100",
		"10000001",
		"10000111",
		"10010000",
		"10010011",
		"10010010",
		"10010011",
		"10010101",
		"10011110",
		"10010011",
		"10000101",
		"01110101",
		"01011101",
		"01010100",
		"01110110",
		"00111100",
		"00100101",
		"01110001",
		"10000110",
		"10001100",
		"10100000",
		"10001100",
		"10000010",
		"10001111",
		"10001100",
		"10001010",
		"10100110",
		"11000010",
		"11000000",
		"11000100",
		"11010001",
		"10010011",
		"10010010",
		"10010111",
		"10000010",
		"01110010",
		"01101110",
		"01101010",
		"01111011",
		"10000111",
		"10010000",
		"10011010",
		"10101000",
		"10101010",
		"10100010",
		"10011000",
		"10010001",
		"10010000",
		"10010111",
		"10011000",
		"10011000",
		"10011000",
		"10011101",
		"10100110",
		"10111100",
		"11001101",
		"11010101",
		"11010100",
		"11010001",
		"11000001",
		"10011010",
		"01111000",
		"00100000",
		"00010100",
		"01000100",
		"01100100",
		"01110011",
		"10000001",
		"10000111",
		"10001001",
		"10001001",
		"10001100",
		"10001111",
		"10001011",
		"10000101",
		"10000001",
		"10000010",
		"10000101",
		"01111110",
		"01110100",
		"01111001",
		"10001101",
		"10011110",
		"10100010",
		"10001010",
		"01011110",
		"01001111",
		"01001111",
		"01010010",
		"01000111",
		"01010010",
		"01101010",
		"01011101",
		"01010010",
		"01001010",
		"01000000",
		"00111001",
		"00110111",
		"00111000",
		"00110111",
		"00111000",
		"00110101",
		"00110110",
		"00111000",
		"00111000",
		"00111001",
		"00111000",
		"00111000",
		"00111010",
		"00111011",
		"00111000",
		"00111000",
		"00110110",
		"00110101",
		"00110000",
		"00101111",
		"10000010",
		"10011101",
		"10101001",
		"10101000",
		"10100110",
		"10100011",
		"10100010",
		"10100010",
		"10100001",
		"10100010",
		"10100101",
		"10100111",
		"10101001",
		"10101101",
		"10101111",
		"10110100",
		"10111000",
		"10111011",
		"10111010",
		"10111011",
		"10111111",
		"10111101",
		"10111100",
		"10111100",
		"10111111",
		"11000001",
		"11000000",
		"10111111",
		"10110001",
		"10001001",
		"00110001",
		"00101101",
		"01000111",
		"01110110",
		"10001010",
		"10001111",
		"10010001",
		"10100000",
		"10100111",
		"10011101",
		"10011100",
		"10011111",
		"10011110",
		"10011011",
		"10011100",
		"10011100",
		"10010000",
		"01011100",
		"00110100",
		"00101111",
		"00111011",
		"01001010",
		"00111100",
		"00101100",
		"01100001",
		"01111111",
		"10001110",
		"10011010",
		"10010011",
		"10001110",
		"10100001",
		"10110101",
		"11001010",
		"11000110",
		"11001111",
		"11000001",
		"10110000",
		"01110001",
		"01001001",
		"10001110",
		"10011011",
		"01111010",
		"01110111",
		"10000110",
		"10010001",
		"10011010",
		"10000110",
		"01101100",
		"01011010",
		"01010111",
		"01011011",
		"01101001",
		"10000110",
		"10010111",
		"10010110",
		"10010010",
		"10010011",
		"10010100",
		"10011100",
		"10110001",
		"11001101",
		"11011001",
		"11011000",
		"11010001",
		"10100111",
		"10001101",
		"00111010",
		"00001001",
		"00100011",
		"01001111",
		"01100011",
		"01110010",
		"01110110",
		"01110101",
		"01110011",
		"01110101",
		"01110100",
		"01101101",
		"01100110",
		"01100110",
		"01100100",
		"01011010",
		"01010001",
		"01011010",
		"01110001",
		"01111001",
		"01101011",
		"01100100",
		"01010100",
		"01001111",
		"01010010",
		"01010010",
		"01010100",
		"01001010",
		"01001011",
		"01010111",
		"01001100",
		"01001000",
		"01000100",
		"01000000",
		"01000000",
		"00111100",
		"00111001",
		"00110110",
		"00110110",
		"00110110",
		"00110111",
		"00110111",
		"00110110",
		"00111010",
		"00111000",
		"00111001",
		"00111011",
		"00111011",
		"00111001",
		"00111001",
		"00110111",
		"00110100",
		"00101110",
		"00110011",
		"10000100",
		"10011101",
		"10101000",
		"10101000",
		"10100101",
		"10100011",
		"10100011",
		"10100011",
		"10100010",
		"10100101",
		"10100110",
		"10101010",
		"10101010",
		"10101100",
		"10101110",
		"10110010",
		"10110110",
		"10111001",
		"10111000",
		"10111010",
		"10111110",
		"10111110",
		"10111100",
		"10111100",
		"11000000",
		"11000001",
		"11000001",
		"10111101",
		"10100001",
		"01001110",
		"00010110",
		"00110110",
		"01110101",
		"10000111",
		"10001111",
		"10010010",
		"10011100",
		"10100111",
		"10100111",
		"10100110",
		"10100110",
		"10100101",
		"10100110",
		"10100111",
		"10101010",
		"10110101",
		"11000000",
		"10001101",
		"00111000",
		"01001111",
		"00111000",
		"00011101",
		"00010001",
		"00110111",
		"10000011",
		"10001001",
		"10010100",
		"10011010",
		"10010111",
		"10011000",
		"10100110",
		"10110010",
		"11000110",
		"11001111",
		"11001110",
		"11001000",
		"10111101",
		"10100001",
		"01101101",
		"10001001",
		"10100101",
		"01111011",
		"01101000",
		"01111011",
		"10010011",
		"10010000",
		"01000001",
		"00111110",
		"01000111",
		"01010001",
		"01100001",
		"01110110",
		"10001000",
		"10010000",
		"10011000",
		"10011101",
		"10011111",
		"10100010",
		"10011111",
		"10011010",
		"10100010",
		"10111110",
		"11011010",
		"11010100",
		"10101000",
		"10011000",
		"01010110",
		"00001000",
		"00001111",
		"00110000",
		"01010000",
		"01011100",
		"01011111",
		"01011101",
		"01011111",
		"01011101",
		"01010111",
		"01010001",
		"01010000",
		"01001110",
		"01001010",
		"01001100",
		"01010110",
		"01011011",
		"01011001",
		"01001011",
		"01000110",
		"01001101",
		"01010000",
		"01010011",
		"01010110",
		"01010101",
		"01010110",
		"01010100",
		"00111110",
		"01001110",
		"01001011",
		"01001000",
		"01000110",
		"01000100",
		"01000101",
		"01000010",
		"00111101",
		"00110111",
		"00110110",
		"00110110",
		"00110110",
		"00110110",
		"00111000",
		"00111100",
		"00111100",
		"00111011",
		"00111001",
		"00111000",
		"00110111",
		"00110110",
		"00110100",
		"00110100",
		"00110000",
		"00111001",
		"10000111",
		"10011101",
		"10100100",
		"10100111",
		"10100011",
		"10100010",
		"10100010",
		"10100010",
		"10100010",
		"10100101",
		"10101010",
		"10101101",
		"10101101",
		"10101110",
		"10110001",
		"10110101",
		"10111000",
		"10111010",
		"10111010",
		"10111100",
		"10111110",
		"10111101",
		"10111100",
		"10111101",
		"10111111",
		"11000000",
		"11000001",
		"10111001",
		"01110101",
		"00011111",
		"00011101",
		"01100111",
		"10000101",
		"10001010",
		"10010010",
		"10010111",
		"10011111",
		"10100001",
		"10100100",
		"10100111",
		"10101010",
		"10101100",
		"10110000",
		"10110001",
		"10110010",
		"10110111",
		"10110000",
		"10000011",
		"10010101",
		"10011010",
		"01010110",
		"00011011",
		"00010110",
		"01101100",
		"10001110",
		"10010101",
		"10010011",
		"10100000",
		"10010110",
		"10011011",
		"10100101",
		"10110101",
		"11000110",
		"11010000",
		"11001101",
		"11001000",
		"11000010",
		"11000011",
		"10100110",
		"01101101",
		"10010101",
		"10010000",
		"10001101",
		"10001101",
		"01111101",
		"01000110",
		"00111100",
		"01001011",
		"01010011",
		"01011110",
		"01110101",
		"10000101",
		"10001110",
		"10011000",
		"10011111",
		"10100011",
		"10101000",
		"10101001",
		"10101001",
		"10100111",
		"10100101",
		"10100010",
		"10110001",
		"11001010",
		"10101010",
		"10011101",
		"01100111",
		"00001100",
		"00001011",
		"00011010",
		"00111010",
		"01001010",
		"01001011",
		"01001100",
		"01010000",
		"01001001",
		"01000011",
		"00111110",
		"00110111",
		"00110111",
		"01000110",
		"01010000",
		"01001110",
		"01001101",
		"01001010",
		"01001010",
		"01001111",
		"01010100",
		"01010101",
		"01010111",
		"01011001",
		"01011001",
		"01011001",
		"01010101",
		"00111000",
		"01001111",
		"01010000",
		"01001110",
		"01001100",
		"01001000",
		"01000110",
		"01000101",
		"01000100",
		"00111111",
		"00111000",
		"00110101",
		"00110110",
		"00110110",
		"00111010",
		"01000000",
		"01000010",
		"00111111",
		"00111000",
		"00110111",
		"00110110",
		"00110101",
		"00110110",
		"00110110",
		"00110101",
		"01000101",
		"10001001",
		"10011110",
		"10100001",
		"10100100",
		"10100100",
		"10100001",
		"10100001",
		"10100001",
		"10100010",
		"10100100",
		"10101010",
		"10101101",
		"10101111",
		"10110001",
		"10110011",
		"10110111",
		"10111011",
		"10111100",
		"10111011",
		"10111101",
		"10111101",
		"10111011",
		"10111100",
		"10111100",
		"10111111",
		"10111111",
		"11000011",
		"10011111",
		"00110100",
		"00001100",
		"01000101",
		"10000011",
		"10001101",
		"10010100",
		"10010111",
		"10011010",
		"10011000",
		"10010100",
		"10010101",
		"10011001",
		"10011100",
		"10100010",
		"10100101",
		"10101010",
		"10100101",
		"10000001",
		"00111000",
		"01011101",
		"10101111",
		"10111101",
		"10011011",
		"01110010",
		"01000111",
		"00111100",
		"01111010",
		"10010100",
		"10101001",
		"10101110",
		"10100011",
		"10100010",
		"10101001",
		"10110001",
		"10111011",
		"11001101",
		"11000111",
		"10111010",
		"10111010",
		"11001000",
		"10111110",
		"01111111",
		"10010000",
		"10100110",
		"10011010",
		"10000110",
		"10001111",
		"01000000",
		"01010001",
		"01011111",
		"01101000",
		"01101110",
		"01110011",
		"10000001",
		"10000111",
		"10010010",
		"10011010",
		"10100010",
		"10100101",
		"10101000",
		"10101011",
		"10101111",
		"10101100",
		"10100110",
		"10100110",
		"10101010",
		"10011110",
		"10011001",
		"01011110",
		"00001001",
		"00001110",
		"00010110",
		"00101011",
		"00111001",
		"00111111",
		"01000010",
		"01000001",
		"00111110",
		"00111000",
		"00101111",
		"00110011",
		"01000000",
		"01000110",
		"01001001",
		"01001001",
		"01001001",
		"01001111",
		"01010010",
		"01010010",
		"01010110",
		"01010101",
		"01010111",
		"01011000",
		"01011011",
		"01011010",
		"01010111",
		"00110011",
		"01001110",
		"01001010",
		"01001100",
		"01001101",
		"01001011",
		"01001010",
		"01000110",
		"01000111",
		"01000110",
		"01000000",
		"00111100",
		"00111000",
		"00111001",
		"00111110",
		"01000101",
		"01000110",
		"01000011",
		"00111001",
		"00110110",
		"00110111",
		"00110111",
		"00111000",
		"00111001",
		"00110011",
		"01000110",
		"10001110",
		"10011110",
		"10100011",
		"10100110",
		"10100101",
		"10100011",
		"10100010",
		"10100100",
		"10100100",
		"10101000",
		"10101100",
		"10101110",
		"10110000",
		"10110011",
		"10110110",
		"10111001",
		"10111100",
		"10111100",
		"10111011",
		"10111101",
		"10111100",
		"10111100",
		"10111101",
		"10111101",
		"11000000",
		"11000000",
		"10111111",
		"01110010",
		"00010001",
		"00010001",
		"01100011",
		"10001111",
		"10010101",
		"10010110",
		"10010110",
		"10010111",
		"10010001",
		"10001110",
		"10001101",
		"10010001",
		"10011010",
		"10011111",
		"10100010",
		"10100101",
		"10101011",
		"10110001",
		"10010010",
		"01000110",
		"00101010",
		"01100011",
		"10011000",
		"10100011",
		"10100011",
		"01111110",
		"10001011",
		"10100101",
		"10100101",
		"10000001",
		"10010001",
		"10100011",
		"10101111",
		"10101111",
		"10111010",
		"11001001",
		"11001010",
		"11000111",
		"10101000",
		"10010100",
		"10000100",
		"10011001",
		"10110001",
		"10111000",
		"10101000",
		"10010000",
		"01011101",
		"01001001",
		"01101101",
		"01110101",
		"01110100",
		"01111001",
		"01111001",
		"10000001",
		"10001100",
		"10010110",
		"10100000",
		"10100010",
		"10100110",
		"10101001",
		"10101010",
		"10101100",
		"10101111",
		"10101110",
		"10100111",
		"10100111",
		"10011111",
		"10001101",
		"01000101",
		"00001000",
		"00001100",
		"00010000",
		"00011011",
		"00101011",
		"00110010",
		"00110101",
		"00110100",
		"00101101",
		"00100110",
		"00101110",
		"00111110",
		"01000001",
		"01000111",
		"01001100",
		"01001110",
		"01010001",
		"01010010",
		"01010100",
		"01010010",
		"01010101",
		"01010100",
		"01010110",
		"01010110",
		"01011001",
		"01011100",
		"01010110",
		"00110000",
		"01001011",
		"01000111",
		"01000000",
		"01000110",
		"01001110",
		"01001101",
		"01001001",
		"01000111",
		"01001010",
		"01001000",
		"01000011",
		"00111011",
		"00111100",
		"00111111",
		"01001001",
		"01001000",
		"00111110",
		"00111000",
		"00111000",
		"00111001",
		"00110111",
		"00110110",
		"00110011",
		"00101011",
		"01010000",
		"10001111",
		"10100000",
		"10101001",
		"10100110",
		"10100010",
		"10100001",
		"10100011",
		"10100101",
		"10100101",
		"10101000",
		"10101011",
		"10110000",
		"10110010",
		"10110101",
		"10111000",
		"10111010",
		"10111011",
		"10111010",
		"10111011",
		"10111110",
		"10111101",
		"10111100",
		"10111101",
		"10111101",
		"10111110",
		"10111101",
		"10101010",
		"01000011",
		"00001000",
		"00110011",
		"01111001",
		"10011001",
		"10011101",
		"10011101",
		"10011110",
		"10011101",
		"10011000",
		"10010110",
		"10010110",
		"10010110",
		"10011000",
		"10011001",
		"10011101",
		"10011111",
		"10100100",
		"10100101",
		"10101110",
		"10101101",
		"01101011",
		"00111000",
		"01010010",
		"01101101",
		"01111100",
		"10000111",
		"01111110",
		"10010010",
		"10101100",
		"10011101",
		"10100001",
		"10110001",
		"10111100",
		"10111110",
		"10110100",
		"10101110",
		"10110110",
		"11000000",
		"10000001",
		"01111110",
		"10010110",
		"10100101",
		"10100110",
		"10000010",
		"10001101",
		"00110011",
		"00000110",
		"00111011",
		"01101000",
		"01101101",
		"01101001",
		"01101010",
		"01111000",
		"10001110",
		"10010100",
		"10011010",
		"10100011",
		"10100111",
		"10101011",
		"10110000",
		"10110011",
		"10110100",
		"10110100",
		"10110010",
		"10101111",
		"10101010",
		"10101000",
		"10000001",
		"00101000",
		"00001000",
		"00001011",
		"00001110",
		"00010011",
		"00011001",
		"00100000",
		"00100101",
		"00100101",
		"00011011",
		"00110000",
		"01000001",
		"01000100",
		"01001001",
		"01001000",
		"01001011",
		"01010001",
		"01010010",
		"01010001",
		"01010100",
		"01010010",
		"01010011",
		"01010011",
		"01010101",
		"01010100",
		"01011000",
		"01011011",
		"01011011",
		"00110011",
		"01000111",
		"01000111",
		"01000100",
		"01000010",
		"01000101",
		"01001001",
		"01001010",
		"01001001",
		"01001011",
		"01001001",
		"01000101",
		"00111101",
		"00111010",
		"00111011",
		"01000100",
		"01000010",
		"00111011",
		"00111000",
		"00110111",
		"00110110",
		"00110100",
		"00101111",
		"00101011",
		"00100011",
		"01100010",
		"10010001",
		"10100000",
		"10101011",
		"10100101",
		"10100001",
		"10100010",
		"10100011",
		"10100100",
		"10100110",
		"10101000",
		"10101011",
		"10110000",
		"10110101",
		"10110110",
		"10111000",
		"10111010",
		"10111001",
		"10111001",
		"10111010",
		"10111101",
		"10111101",
		"10111101",
		"10111011",
		"10111011",
		"10111010",
		"10101110",
		"10000011",
		"00011110",
		"00010111",
		"01101110",
		"10010000",
		"10011110",
		"10100000",
		"10100001",
		"10100000",
		"10011100",
		"10010101",
		"10010100",
		"10010110",
		"10010110",
		"10010101",
		"10010000",
		"10001001",
		"10000010",
		"01111111",
		"01111111",
		"01111101",
		"10000111",
		"10011011",
		"10011111",
		"10011101",
		"10011110",
		"10011010",
		"10010001",
		"10000011",
		"10001011",
		"10011100",
		"10100001",
		"10011111",
		"10011000",
		"10000001",
		"01111011",
		"01100110",
		"10000010",
		"10011001",
		"10010101",
		"10000000",
		"10001000",
		"10011010",
		"10010101",
		"10000101",
		"01111100",
		"10010000",
		"10001101",
		"01101101",
		"01101110",
		"01111100",
		"10000111",
		"10001101",
		"10001101",
		"10010001",
		"10010100",
		"10011000",
		"10011011",
		"10011111",
		"10100100",
		"10101011",
		"10110010",
		"10111001",
		"11000000",
		"11000001",
		"10111011",
		"10110010",
		"10101100",
		"10101010",
		"10001110",
		"00011100",
		"00001001",
		"00001100",
		"00001101",
		"00001111",
		"00010001",
		"00010011",
		"00010011",
		"00010010",
		"00110000",
		"01001100",
		"01001011",
		"01001001",
		"01001000",
		"01001001",
		"01001101",
		"01010000",
		"01010010",
		"01010100",
		"01010101",
		"01010100",
		"01010100",
		"01010101",
		"01010110",
		"01010101",
		"01010111",
		"01100011",
		"01101110",
		"00110100",
		"01000010",
		"00111110",
		"01000011",
		"00111111",
		"01000000",
		"01000010",
		"01000100",
		"01000101",
		"01000111",
		"01001000",
		"01000100",
		"00111101",
		"00111001",
		"00111001",
		"00111101",
		"00111111",
		"00111001",
		"00111000",
		"00110101",
		"00110001",
		"00101111",
		"00101001",
		"00100101",
		"00100000",
		"01101110",
		"10010010",
		"10100101",
		"10101011",
		"10100110",
		"10100010",
		"10100011",
		"10100101",
		"10100011",
		"10100110",
		"10101010",
		"10101101",
		"10110001",
		"10110101",
		"10111000",
		"10111010",
		"10111010",
		"10111001",
		"10111011",
		"10111101",
		"10111101",
		"10111011",
		"10111010",
		"10111001",
		"10110111",
		"10101111",
		"10010110",
		"01001111",
		"00001011",
		"00110100",
		"10000000",
		"10011100",
		"10100111",
		"10100000",
		"10011011",
		"10010100",
		"10001101",
		"10001111",
		"10010001",
		"10010011",
		"10010110",
		"10010101",
		"10001111",
		"10001110",
		"10001011",
		"10001001",
		"10001011",
		"10001110",
		"10010010",
		"10010011",
		"10010111",
		"10011000",
		"10011000",
		"10010100",
		"10010001",
		"10010100",
		"10011001",
		"10011001",
		"10011011",
		"10011100",
		"10100101",
		"10100110",
		"10001001",
		"00110001",
		"00001000",
		"00110111",
		"01101001",
		"01101011",
		"01101110",
		"01110101",
		"10000100",
		"10010011",
		"10011010",
		"10100001",
		"10011110",
		"10100010",
		"10100100",
		"10100001",
		"10011111",
		"10100010",
		"10100001",
		"10100000",
		"10011110",
		"10011111",
		"10100001",
		"10100000",
		"10100100",
		"10101110",
		"10110100",
		"10110110",
		"11000011",
		"11001000",
		"11000010",
		"10110101",
		"10101100",
		"10101001",
		"10011110",
		"00100111",
		"00000111",
		"00001010",
		"00001011",
		"00001101",
		"00001100",
		"00001100",
		"00001101",
		"00110011",
		"01010011",
		"01001001",
		"01001001",
		"01001011",
		"01001110",
		"01001111",
		"01001111",
		"01010001",
		"01010110",
		"01010111",
		"01010110",
		"01011000",
		"01010111",
		"01010111",
		"01010110",
		"01010111",
		"01011100",
		"01111001",
		"10010000",
		"00111000",
		"01000010",
		"00111010",
		"00111010",
		"00111001",
		"00111101",
		"00111100",
		"00111110",
		"01000011",
		"01000100",
		"01000011",
		"01000000",
		"00111111",
		"00111100",
		"00111010",
		"00111001",
		"00111011",
		"00111010",
		"00110111",
		"00110011",
		"00101110",
		"00101101",
		"00100111",
		"00100101",
		"00100101",
		"01111010",
		"10010011",
		"10101010",
		"10101010",
		"10100101",
		"10100011",
		"10100011",
		"10100100",
		"10100011",
		"10100110",
		"10101011",
		"10101111",
		"10110001",
		"10110110",
		"10111001",
		"10111010",
		"10111010",
		"10111001",
		"10111011",
		"10111101",
		"10111100",
		"10111011",
		"10111001",
		"10110111",
		"10101111",
		"10011110",
		"01110101",
		"00101000",
		"00001111",
		"01010010",
		"10000110",
		"10011111",
		"10101000",
		"10011100",
		"10001110",
		"10001000",
		"10001101",
		"10001100",
		"10010010",
		"10010101",
		"10010001",
		"10010001",
		"10010000",
		"10001101",
		"10001100",
		"10001101",
		"10001101",
		"10010000",
		"10010000",
		"10001111",
		"10010110",
		"10010110",
		"10010111",
		"10011010",
		"10011101",
		"10011111",
		"10011101",
		"10011101",
		"10011011",
		"10011110",
		"10100010",
		"10100101",
		"10101100",
		"10100011",
		"01110100",
		"01010001",
		"01101110",
		"01110111",
		"01111000",
		"01111110",
		"10000101",
		"10001111",
		"10011000",
		"10100000",
		"10100011",
		"10100001",
		"10100001",
		"10100110",
		"10100100",
		"10100010",
		"10100011",
		"10100111",
		"10100110",
		"10100101",
		"10100100",
		"10100010",
		"10100100",
		"10100111",
		"10110010",
		"10111000",
		"11000001",
		"11000100",
		"11000011",
		"10110100",
		"10110010",
		"10101011",
		"10100010",
		"01000000",
		"00000101",
		"00001010",
		"00001011",
		"00001011",
		"00001010",
		"00001010",
		"00110000",
		"01010000",
		"01001000",
		"01000110",
		"01001000",
		"01001100",
		"01001111",
		"01010000",
		"01010010",
		"01010010",
		"01010011",
		"01011000",
		"01011101",
		"01011011",
		"01011011",
		"01011010",
		"01011100",
		"01100001",
		"10000011",
		"10110000",
		"10111011",
		"00111001",
		"01000010",
		"00111010",
		"00111001",
		"00111100",
		"00111110",
		"00111010",
		"00111011",
		"01000000",
		"01000010",
		"01000001",
		"00111111",
		"00111110",
		"00111100",
		"00111010",
		"00111010",
		"00111000",
		"00111000",
		"00110111",
		"00110001",
		"00101101",
		"00101001",
		"00100111",
		"00011110",
		"00101110",
		"10000011",
		"10010101",
		"10101010",
		"10101001",
		"10100011",
		"10100010",
		"10100010",
		"10100011",
		"10100101",
		"10101000",
		"10101100",
		"10101111",
		"10110010",
		"10110110",
		"10111000",
		"10111010",
		"10111000",
		"10110111",
		"10111001",
		"10111011",
		"10111011",
		"10111001",
		"10110110",
		"10110001",
		"10100001",
		"10001000",
		"01010001",
		"00010111",
		"00011110",
		"01100110",
		"10001000",
		"10011000",
		"10011011",
		"10001110",
		"10001001",
		"10001010",
		"10001011",
		"10001100",
		"10001111",
		"10001110",
		"10001101",
		"10001010",
		"10000100",
		"10000101",
		"10001010",
		"10001001",
		"10001100",
		"10001100",
		"10001011",
		"10010000",
		"10010100",
		"10010010",
		"10010011",
		"10011001",
		"10011111",
		"10011101",
		"10011011",
		"10011011",
		"10011111",
		"10100111",
		"10110011",
		"10110101",
		"10101110",
		"10101000",
		"10010110",
		"01100001",
		"01101010",
		"01110101",
		"01111100",
		"10000010",
		"10001011",
		"10001101",
		"10010011",
		"10011001",
		"10100010",
		"10100110",
		"10100111",
		"10101001",
		"10101111",
		"10110010",
		"10110011",
		"10110111",
		"10111110",
		"11000000",
		"10111111",
		"10111111",
		"10110100",
		"10101010",
		"10101110",
		"10110101",
		"11000000",
		"11000001",
		"11000001",
		"10110111",
		"10111010",
		"10110010",
		"10100100",
		"01010001",
		"00000110",
		"00001010",
		"00001011",
		"00001011",
		"00001100",
		"00110000",
		"01001000",
		"01000000",
		"00111111",
		"01000010",
		"01000111",
		"01001100",
		"01010000",
		"01010000",
		"01010001",
		"01010101",
		"01010100",
		"01010110",
		"01011010",
		"01011100",
		"01011101",
		"01011100",
		"01100100",
		"10000001",
		"10111010",
		"11010010",
		"11010010",
		"00110100",
		"01000100",
		"00111100",
		"00111100",
		"01000001",
		"00111010",
		"00110110",
		"00110011",
		"00110010",
		"00111101",
		"01000000",
		"00111110",
		"00111100",
		"00111010",
		"00111010",
		"00110110",
		"00110101",
		"00110100",
		"00110011",
		"00101111",
		"00101011",
		"00100101",
		"00100110",
		"00011010",
		"01000011",
		"10001011",
		"10010111",
		"10101000",
		"10100110",
		"10100010",
		"10100010",
		"10100010",
		"10100011",
		"10100110",
		"10101010",
		"10101110",
		"10110000",
		"10110100",
		"10110110",
		"10111000",
		"10111001",
		"10110110",
		"10110110",
		"10111001",
		"10111010",
		"10111000",
		"10110101",
		"10110000",
		"10100101",
		"10010001",
		"01101110",
		"00110111",
		"00010001",
		"00110000",
		"01110000",
		"10000010",
		"10001100",
		"10001000",
		"10000011",
		"10001000",
		"10001000",
		"10001010",
		"10001100",
		"10001001",
		"10001011",
		"10001010",
		"10001000",
		"10000111",
		"10001001",
		"10001100",
		"10001110",
		"10001110",
		"10001111",
		"10010100",
		"10010111",
		"10010101",
		"10001111",
		"10010101",
		"10011001",
		"10011101",
		"10011001",
		"10011001",
		"10011101",
		"10100010",
		"10111001",
		"11010000",
		"11010101",
		"11001110",
		"11000101",
		"10110000",
		"01110111",
		"01100100",
		"01110010",
		"01111011",
		"10000101",
		"10001011",
		"10001010",
		"10001101",
		"10010111",
		"10011110",
		"10100100",
		"10100111",
		"10101000",
		"10111001",
		"11001001",
		"11010101",
		"11010111",
		"11011000",
		"11011000",
		"11011000",
		"11010101",
		"11001010",
		"10110100",
		"10101110",
		"10110001",
		"10111101",
		"10111110",
		"10111011",
		"10110110",
		"10110101",
		"10101111",
		"10100010",
		"01011001",
		"00001000",
		"00001011",
		"00001010",
		"00001110",
		"00110001",
		"01000110",
		"00111100",
		"00111101",
		"00111111",
		"01000010",
		"01000110",
		"01001011",
		"01010011",
		"01010101",
		"01010110",
		"01010100",
		"01010101",
		"01011001",
		"01011001",
		"01011100",
		"01011101",
		"01101001",
		"01111000",
		"10100110",
		"11001010",
		"11011010",
		"11010101",
		"00110100",
		"01000100",
		"00111101",
		"00111111",
		"00111111",
		"00111100",
		"00111010",
		"00110011",
		"00101001",
		"00100111",
		"00111001",
		"00111110",
		"00111100",
		"00111010",
		"00111000",
		"00110010",
		"00101010",
		"00100001",
		"00100001",
		"00100100",
		"00100001",
		"00011011",
		"00011100",
		"00010011",
		"01011101",
		"10001100",
		"10011000",
		"10100111",
		"10101000",
		"10100011",
		"10100011",
		"10100011",
		"10100101",
		"10100111",
		"10101011",
		"10101101",
		"10110000",
		"10110100",
		"10110111",
		"10111001",
		"10111001",
		"10110111",
		"10111000",
		"10111100",
		"10110110",
		"10110101",
		"10110001",
		"10100111",
		"10010110",
		"01111111",
		"01010101",
		"00100011",
		"00010001",
		"00111111",
		"01110000",
		"01111101",
		"10000010",
		"10000011",
		"10000110",
		"10001010",
		"10001100",
		"10001010",
		"10001000",
		"10001011",
		"10001011",
		"10001001",
		"10000111",
		"10001010",
		"10001011",
		"10001100",
		"10001101",
		"10001110",
		"10010000",
		"10010110",
		"10010111",
		"10010110",
		"10010100",
		"10010110",
		"10011000",
		"10010100",
		"10010111",
		"10011100",
		"10100001",
		"10101010",
		"11000001",
		"11010110",
		"11011010",
		"11011010",
		"11011000",
		"11010101",
		"10010010",
		"01100011",
		"01110110",
		"01111101",
		"10000011",
		"10000000",
		"10000001",
		"10000111",
		"10010001",
		"10011001",
		"10100010",
		"10100111",
		"10101010",
		"10110010",
		"11000011",
		"11010101",
		"11011011",
		"11011001",
		"11010111",
		"11010100",
		"11001111",
		"11000011",
		"10110000",
		"10101001",
		"10101101",
		"10110101",
		"10111100",
		"10110100",
		"10101110",
		"10110000",
		"10100110",
		"10100010",
		"01011000",
		"00001010",
		"00001110",
		"00001110",
		"00101100",
		"00111111",
		"00111010",
		"00111011",
		"00111100",
		"00111110",
		"01000010",
		"01000111",
		"01001100",
		"01010011",
		"01011000",
		"01011000",
		"01010110",
		"01010110",
		"01011001",
		"01011010",
		"01011010",
		"01011110",
		"01110111",
		"10100110",
		"10111100",
		"11010100",
		"11011100",
		"11001100",
		"00111010",
		"01000101",
		"00111110",
		"00111101",
		"00111111",
		"01000001",
		"01000100",
		"00111011",
		"00101111",
		"00100101",
		"00100000",
		"00101101",
		"00110110",
		"00110101",
		"00110000",
		"00100110",
		"00100110",
		"00101010",
		"00110010",
		"00111110",
		"01001111",
		"01001111",
		"00101101",
		"00001110",
		"01101111",
		"10001011",
		"10011001",
		"10100101",
		"10101000",
		"10100011",
		"10100101",
		"10100101",
		"10100111",
		"10101001",
		"10101101",
		"10101100",
		"10101111",
		"10110011",
		"10110110",
		"10110111",
		"10110111",
		"10110110",
		"10110111",
		"10110110",
		"10110010",
		"10101111",
		"10101000",
		"10011001",
		"10001010",
		"01110001",
		"01000110",
		"00011011",
		"00010101",
		"01001010",
		"01110000",
		"01111001",
		"01111101",
		"10000100",
		"10001010",
		"10001001",
		"10001001",
		"10001011",
		"10001101",
		"10001110",
		"10001010",
		"10000111",
		"10001011",
		"10001010",
		"10000111",
		"10001001",
		"10001010",
		"10001101",
		"10010001",
		"10010101",
		"10010111",
		"10010100",
		"10010011",
		"10010101",
		"10010110",
		"10010010",
		"10011000",
		"10100010",
		"10110010",
		"10111011",
		"11000101",
		"11010001",
		"11010110",
		"11010110",
		"11011001",
		"11011001",
		"10100110",
		"01011110",
		"01110001",
		"01111001",
		"01110110",
		"01111000",
		"01111101",
		"10000100",
		"10001010",
		"10010000",
		"10011001",
		"10100010",
		"10101001",
		"10110000",
		"10111011",
		"11000110",
		"11001100",
		"11001101",
		"11001011",
		"11000011",
		"10110110",
		"10101110",
		"10100111",
		"10100111",
		"10101011",
		"10101110",
		"10110101",
		"10110000",
		"10101111",
		"10101100",
		"10100100",
		"10100011",
		"01010001",
		"00001011",
		"00001111",
		"00011111",
		"00111001",
		"00111000",
		"00111010",
		"00111101",
		"01000010",
		"01000101",
		"01000111",
		"01001011",
		"01001110",
		"01010101",
		"01011011",
		"01011010",
		"01011001",
		"01011001",
		"01011011",
		"01011101",
		"01011110",
		"01100011",
		"01111100",
		"10110010",
		"11001100",
		"11011000",
		"11010101",
		"10101100",
		"00111011",
		"01000101",
		"00111110",
		"00111101",
		"00111101",
		"01000001",
		"01000111",
		"00111111",
		"00110011",
		"00101001",
		"00011100",
		"00010001",
		"00100100",
		"00111101",
		"01001101",
		"01001100",
		"00111100",
		"00111110",
		"01010001",
		"01011001",
		"01001101",
		"00101100",
		"00010100",
		"00100000",
		"10000011",
		"10001011",
		"10011010",
		"10100100",
		"10100100",
		"10100001",
		"10100100",
		"10100100",
		"10100111",
		"10101010",
		"10101100",
		"10101101",
		"10110000",
		"10110011",
		"10110100",
		"10110101",
		"10110011",
		"10110000",
		"10110010",
		"10110010",
		"10101111",
		"10101010",
		"10100000",
		"10010011",
		"10000001",
		"01101000",
		"01000001",
		"00011001",
		"00011100",
		"01001100",
		"01101101",
		"01111000",
		"01111110",
		"10001000",
		"10001011",
		"10001011",
		"10001100",
		"10001111",
		"10010000",
		"10001101",
		"10000111",
		"10000111",
		"10001000",
		"10001001",
		"10001000",
		"10001010",
		"10001101",
		"10010001",
		"10010000",
		"10010011",
		"10010010",
		"10001110",
		"10001011",
		"10010000",
		"10010101",
		"10011011",
		"10011111",
		"10101011",
		"10111001",
		"10111010",
		"10111100",
		"10111011",
		"11000000",
		"11000101",
		"11001100",
		"11001101",
		"10110001",
		"01110001",
		"01100110",
		"01110000",
		"01101111",
		"01110010",
		"01110111",
		"01111010",
		"10000001",
		"10000111",
		"10010001",
		"10010101",
		"10010110",
		"10011010",
		"10100110",
		"10101001",
		"10110000",
		"10110110",
		"10110100",
		"10101101",
		"10101000",
		"10101000",
		"10101011",
		"10100111",
		"10100101",
		"10101001",
		"10101100",
		"10101100",
		"10101010",
		"10100111",
		"10100100",
		"10100011",
		"01000100",
		"00000111",
		"00001101",
		"00101001",
		"00110001",
		"00110000",
		"00111000",
		"00111101",
		"01000011",
		"01001001",
		"01001100",
		"01001110",
		"01010000",
		"01010101",
		"01011011",
		"01011011",
		"01011010",
		"01011000",
		"01011100",
		"01100001",
		"01100011",
		"01101111",
		"10010001",
		"10111000",
		"11000111",
		"11000111",
		"10101100",
		"01110000",
		"00111101",
		"01000011",
		"01000001",
		"00111110",
		"00111100",
		"00111100",
		"00111110",
		"00111001",
		"00110001",
		"00100001",
		"00100101",
		"00111100",
		"01001000",
		"00111101",
		"00111011",
		"01000111",
		"00111011",
		"00100110",
		"00110001",
		"01001111",
		"00101110",
		"00010101",
		"00001110",
		"00111000",
		"10001011",
		"10001110",
		"10011110",
		"10100100",
		"10100110",
		"10100100",
		"10100101",
		"10100100",
		"10101000",
		"10101100",
		"10101101",
		"10101101",
		"10110001",
		"10110100",
		"10110100",
		"10110011",
		"10101111",
		"10101101",
		"10101111",
		"10110001",
		"10101100",
		"10100011",
		"10011010",
		"10001110",
		"01111110",
		"01100100",
		"00111110",
		"00010101",
		"00011111",
		"01001110",
		"01101100",
		"01110100",
		"01111011",
		"10000100",
		"10001101",
		"10001101",
		"10001111",
		"10010010",
		"10010000",
		"10001110",
		"10001100",
		"10001001",
		"10001001",
		"10000111",
		"10000111",
		"10001000",
		"10001011",
		"10001111",
		"10010000",
		"10010000",
		"10001100",
		"10000100",
		"10001000",
		"10001111",
		"10010101",
		"10011011",
		"10011111",
		"10100101",
		"10100011",
		"10101000",
		"10101000",
		"10100111",
		"10101010",
		"10110011",
		"10110111",
		"10110110",
		"10101110",
		"01111101",
		"01100010",
		"01101010",
		"01101010",
		"01101101",
		"01110100",
		"01110101",
		"01111011",
		"10000101",
		"10001011",
		"10001100",
		"10010000",
		"10001111",
		"10010011",
		"10010111",
		"10011010",
		"10100010",
		"10100110",
		"10101000",
		"10100111",
		"10100110",
		"10100111",
		"10100101",
		"10100100",
		"10100110",
		"10100110",
		"10100101",
		"10100011",
		"10100100",
		"10100011",
		"10011101",
		"00101110",
		"00000110",
		"00010000",
		"00101001",
		"00101010",
		"00101111",
		"00110100",
		"00111100",
		"01000011",
		"01001010",
		"01001101",
		"01001110",
		"01010001",
		"01010111",
		"01011010",
		"01011011",
		"01011010",
		"01011010",
		"01011110",
		"01100010",
		"01100111",
		"10000010",
		"10101011",
		"10111001",
		"10111111",
		"10100101",
		"01110011",
		"01011010",
		"00111000",
		"01000000",
		"00111111",
		"01000000",
		"00111111",
		"00111110",
		"00111000",
		"00110100",
		"00100111",
		"00111010",
		"01100111",
		"01010010",
		"00100111",
		"00100110",
		"01010100",
		"01101001",
		"01100100",
		"01001010",
		"01011011",
		"01101110",
		"01000000",
		"00010111",
		"00010010",
		"01010011",
		"10010000",
		"10010011",
		"10100001",
		"10100101",
		"10100101",
		"10100101",
		"10100110",
		"10100100",
		"10101000",
		"10101100",
		"10101101",
		"10101110",
		"10110010",
		"10110010",
		"10110010",
		"10110010",
		"10101101",
		"10101011",
		"10101101",
		"10101101",
		"10100111",
		"10011110",
		"10010101",
		"10001010",
		"01111100",
		"01100100",
		"00111100",
		"00010111",
		"00100000",
		"01001101",
		"01100111",
		"01110010",
		"01111001",
		"01111001",
		"10000011",
		"10000101",
		"10000110",
		"10001011",
		"10001110",
		"10001101",
		"10001101",
		"10001010",
		"10001001",
		"10000111",
		"10000101",
		"10000110",
		"10001001",
		"10000111",
		"10001000",
		"10001011",
		"10000011",
		"01111101",
		"10000111",
		"10010000",
		"10010011",
		"10010101",
		"10011000",
		"10011011",
		"10011001",
		"10011100",
		"10011101",
		"10100001",
		"10100000",
		"10100011",
		"10100100",
		"10100010",
		"10011011",
		"01111111",
		"01101000",
		"01100011",
		"01101000",
		"01101100",
		"01110100",
		"01110111",
		"01111011",
		"10000010",
		"10000101",
		"10001000",
		"10001101",
		"10001100",
		"10001111",
		"10010001",
		"10011000",
		"10011110",
		"10100011",
		"10100101",
		"10100100",
		"10100100",
		"10100100",
		"10100010",
		"10011111",
		"10100001",
		"10100100",
		"10100001",
		"10100000",
		"10100011",
		"10100010",
		"10010110",
		"00100001",
		"00001000",
		"00011001",
		"00100111",
		"00101000",
		"00110001",
		"00111000",
		"01000000",
		"01000100",
		"01001001",
		"01001010",
		"01001110",
		"01010101",
		"01011011",
		"01011010",
		"01011000",
		"01011001",
		"01011100",
		"01011110",
		"01100100",
		"01110010",
		"10010010",
		"10101110",
		"10110001",
		"10100011",
		"01111000",
		"01011111",
		"01011001",
		"00101111",
		"00111100",
		"00111011",
		"00111010",
		"00111000",
		"00111000",
		"00110100",
		"00101100",
		"00111001",
		"01010001",
		"00110111",
		"00010111",
		"00100111",
		"01101101",
		"01011001",
		"01001100",
		"01010101",
		"00100101",
		"00110011",
		"00110111",
		"00100001",
		"00011011",
		"00011101",
		"01100110",
		"10001111",
		"10011000",
		"10100101",
		"10100111",
		"10100111",
		"10100110",
		"10100100",
		"10100111",
		"10101011",
		"10101101",
		"10101110",
		"10110000",
		"10110001",
		"10110001",
		"10110011",
		"10101111",
		"10101011",
		"10101001",
		"10101011",
		"10101010",
		"10100010",
		"10011001",
		"10010001",
		"10001010",
		"01111100",
		"01100001",
		"00110010",
		"00010010",
		"00011100",
		"01000111",
		"01100011",
		"01101111",
		"01110001",
		"01110011",
		"01110101",
		"01110100",
		"01111000",
		"01111010",
		"10000011",
		"10001000",
		"10000110",
		"10000111",
		"10001001",
		"10000101",
		"10000100",
		"10000100",
		"10000011",
		"10000110",
		"10000110",
		"10000101",
		"01111101",
		"01111011",
		"10000000",
		"10001010",
		"10010000",
		"10010001",
		"10010100",
		"10010111",
		"10010110",
		"10010111",
		"10010110",
		"10010111",
		"10010111",
		"10011001",
		"10011011",
		"10010111",
		"10001001",
		"01111001",
		"01101100",
		"01100111",
		"01101010",
		"01110001",
		"01110111",
		"01110101",
		"01111000",
		"01111101",
		"10000010",
		"10000101",
		"10000101",
		"10001001",
		"10001101",
		"10010010",
		"10010111",
		"10011110",
		"10100001",
		"10100010",
		"10100000",
		"10100001",
		"10100001",
		"10011101",
		"10011010",
		"10011010",
		"10100001",
		"10100001",
		"10100001",
		"10100011",
		"10100001",
		"10000101",
		"00010110",
		"00001010",
		"00011011",
		"00100110",
		"00101100",
		"00110100",
		"00111000",
		"01000000",
		"01000010",
		"01000110",
		"01001011",
		"01001111",
		"01010110",
		"01011000",
		"01011001",
		"01011000",
		"01011001",
		"01011011",
		"01011110",
		"01100101",
		"01111001",
		"10011100",
		"10100101",
		"10011011",
		"10000110",
		"01100101",
		"01011100",
		"01010110",
		"00101110",
		"00111001",
		"00110111",
		"00110100",
		"00110000",
		"00101110",
		"00101100",
		"00111111",
		"01011011",
		"00111101",
		"00100101",
		"00011010",
		"01010111",
		"01011110",
		"00100010",
		"01101111",
		"10000010",
		"01100010",
		"01011011",
		"00111111",
		"00011110",
		"00101111",
		"00010011",
		"01110011",
		"10010000",
		"10011001",
		"10101001",
		"10101000",
		"10100110",
		"10100110",
		"10100100",
		"10100110",
		"10101101",
		"10101110",
		"10101110",
		"10110000",
		"10110001",
		"10110010",
		"10110010",
		"10101111",
		"10100111",
		"10100101",
		"10101000",
		"10100111",
		"10011110",
		"10010101",
		"10001101",
		"10000110",
		"01111010",
		"01011111",
		"00101001",
		"00010001",
		"00010011",
		"00110110",
		"01011100",
		"01101101",
		"01101110",
		"01110001",
		"01110000",
		"01101100",
		"01101001",
		"01101010",
		"01110001",
		"01110111",
		"01111011",
		"01111011",
		"01111011",
		"01111001",
		"01111001",
		"01111100",
		"01111100",
		"01111011",
		"01111010",
		"01111010",
		"01111010",
		"01111101",
		"01111101",
		"10000011",
		"10001001",
		"10010000",
		"10010000",
		"10010101",
		"10010111",
		"10010011",
		"10010001",
		"10010001",
		"10001111",
		"10010011",
		"10010001",
		"10001111",
		"10000100",
		"01111001",
		"01101111",
		"01101010",
		"01101010",
		"01101111",
		"01110101",
		"01110011",
		"01110011",
		"01111010",
		"01111111",
		"10000010",
		"10000011",
		"10000111",
		"10001001",
		"10001101",
		"10010010",
		"10010110",
		"10011000",
		"10011011",
		"10011100",
		"10100000",
		"10011110",
		"10011101",
		"10010111",
		"10011010",
		"10100000",
		"10100000",
		"10011111",
		"10100000",
		"10011110",
		"01101101",
		"00010010",
		"00010000",
		"00011011",
		"00101001",
		"00101110",
		"00110101",
		"00111011",
		"01000001",
		"01000010",
		"01000110",
		"01001100",
		"01010010",
		"01010110",
		"01010110",
		"01010111",
		"01011000",
		"01011010",
		"01011101",
		"01011111",
		"01100011",
		"01111010",
		"10011001",
		"10011110",
		"10011111",
		"10000010",
		"01100010",
		"01011001",
		"01010011",
		"00111010",
		"01001011",
		"01000001",
		"00111010",
		"00110110",
		"00110110",
		"00110100",
		"00111110",
		"00110001",
		"00011110",
		"00010100",
		"00101110",
		"01111001",
		"01100010",
		"00111111",
		"01100010",
		"01110011",
		"01111101",
		"01101011",
		"01010010",
		"01000011",
		"00011111",
		"00100100",
		"10000010",
		"10001110",
		"10011011",
		"10101000",
		"10100111",
		"10100101",
		"10100101",
		"10100101",
		"10101000",
		"10101100",
		"10101101",
		"10101110",
		"10110000",
		"10110000",
		"10110001",
		"10101111",
		"10101011",
		"10100111",
		"10101001",
		"10101010",
		"10100100",
		"10011101",
		"10010101",
		"10010000",
		"10001001",
		"01111111",
		"01100010",
		"00101000",
		"00010101",
		"00010010",
		"00101001",
		"01010001",
		"01100110",
		"01101101",
		"01110001",
		"01101010",
		"01100101",
		"01100000",
		"01100010",
		"01100011",
		"01101010",
		"01110010",
		"01110011",
		"01101101",
		"01101110",
		"01101101",
		"01110000",
		"01110001",
		"01110010",
		"01110011",
		"01110010",
		"01110110",
		"01111000",
		"01111101",
		"01111110",
		"10000100",
		"10001100",
		"10010001",
		"10010100",
		"10010111",
		"10010011",
		"10001110",
		"10001110",
		"10001111",
		"10010010",
		"10010000",
		"10001010",
		"10000010",
		"01111011",
		"01110110",
		"01110000",
		"01110010",
		"01111100",
		"01111011",
		"01110110",
		"01110101",
		"01111101",
		"01111111",
		"01111111",
		"10000010",
		"10000111",
		"10001001",
		"10001101",
		"10010001",
		"10010101",
		"10010011",
		"10010100",
		"10011000",
		"10011100",
		"10011110",
		"10011001",
		"10010110",
		"10011010",
		"10011111",
		"10011110",
		"10011101",
		"10011100",
		"10011101",
		"01000111",
		"00001101",
		"00010011",
		"00011010",
		"00100111",
		"00110000",
		"00111000",
		"00111011",
		"00111110",
		"01000100",
		"01001000",
		"01001011",
		"01010001",
		"01010101",
		"01010110",
		"01010110",
		"01010110",
		"01011001",
		"01011101",
		"01100010",
		"01100010",
		"01110010",
		"10001101",
		"10010110",
		"10000101",
		"01100110",
		"01011010",
		"01010100",
		"01010010",
		"00110110",
		"01000011",
		"00111111",
		"00111100",
		"00111100",
		"00111011",
		"00111001",
		"00110001",
		"00111010",
		"00101000",
		"00010111",
		"00110011",
		"01010100",
		"01001001",
		"01000001",
		"01001001",
		"01110001",
		"01111001",
		"01100110",
		"01110101",
		"01100011",
		"00100100",
		"00110100",
		"10001011",
		"10010000",
		"10011100",
		"10101000",
		"10100101",
		"10100100",
		"10100010",
		"10100100",
		"10101000",
		"10101110",
		"10101110",
		"10101111",
		"10110001",
		"10110000",
		"10110001",
		"10101110",
		"10100110",
		"10100110",
		"10101011",
		"10101001",
		"10100100",
		"10011101",
		"10010101",
		"10010001",
		"10001011",
		"10000000",
		"01100000",
		"00100011",
		"00010101",
		"00010010",
		"00011101",
		"01000101",
		"01100000",
		"01101111",
		"01110010",
		"01101111",
		"01100111",
		"01100100",
		"01011110",
		"01011110",
		"01100100",
		"01101100",
		"01101010",
		"01100100",
		"01100111",
		"01100111",
		"01100111",
		"01101101",
		"01110000",
		"01110010",
		"01110010",
		"01110010",
		"01110110",
		"01111000",
		"01111101",
		"10000001",
		"10001011",
		"10010001",
		"10010010",
		"10010001",
		"10001111",
		"10001011",
		"10001011",
		"10001101",
		"10001111",
		"10001101",
		"10000100",
		"01111100",
		"01111000",
		"01110110",
		"01110110",
		"01110101",
		"01111100",
		"01111000",
		"01110111",
		"01111001",
		"01111010",
		"01111111",
		"01111110",
		"10000001",
		"10000110",
		"10001000",
		"10001010",
		"10001101",
		"10010001",
		"10010000",
		"10010011",
		"10010101",
		"10011000",
		"10011001",
		"10010110",
		"10010111",
		"10011000",
		"10011010",
		"10011010",
		"10011100",
		"10011010",
		"10011000",
		"00101110",
		"00001011",
		"00010010",
		"00010111",
		"00101100",
		"00110110",
		"00111010",
		"00111110",
		"00111111",
		"01000100",
		"01001001",
		"01001011",
		"01010000",
		"01010011",
		"01010100",
		"01010101",
		"01010101",
		"01011000",
		"01011010",
		"01011111",
		"01100001",
		"01101100",
		"01111111",
		"01111010",
		"01100111",
		"01011010",
		"01010101",
		"01010001",
		"01001100",
		"00101100",
		"00110011",
		"00110111",
		"00111000",
		"00111000",
		"00110111",
		"00110010",
		"00101010",
		"00101001",
		"00110010",
		"00100101",
		"00100100",
		"00111110",
		"00101010",
		"01001101",
		"01100000",
		"01101111",
		"01110110",
		"01111110",
		"01110101",
		"01011000",
		"01010100",
		"01001100",
		"10001110",
		"10001111",
		"10011010",
		"10101001",
		"10100101",
		"10100101",
		"10100011",
		"10100101",
		"10101010",
		"10101110",
		"10101111",
		"10110000",
		"10101111",
		"10110001",
		"10101111",
		"10101001",
		"10100011",
		"10100100",
		"10100110",
		"10100110",
		"10100011",
		"10011101",
		"10010101",
		"10010001",
		"10001011",
		"10000010",
		"01011000",
		"00011101",
		"00010011",
		"00010010",
		"00010100",
		"00110001",
		"01010010",
		"01100111",
		"01110000",
		"01110001",
		"01101101",
		"01101010",
		"01100100",
		"01011111",
		"01100110",
		"01110001",
		"01101111",
		"01101010",
		"01100100",
		"01100000",
		"01100101",
		"01101011",
		"01110010",
		"01110101",
		"01110010",
		"01110001",
		"01110110",
		"01110101",
		"01111010",
		"10000000",
		"10000101",
		"10001010",
		"10010010",
		"10010010",
		"10010000",
		"10010000",
		"10010010",
		"10001111",
		"10001101",
		"10001001",
		"01111110",
		"01110100",
		"01110001",
		"01110010",
		"01110100",
		"01110111",
		"01111101",
		"01111101",
		"01111001",
		"01111101",
		"01111101",
		"10000001",
		"01111100",
		"01111110",
		"10000101",
		"10001011",
		"10001010",
		"10001110",
		"10010000",
		"10010000",
		"10001111",
		"10010011",
		"10010101",
		"10010111",
		"10010111",
		"10010110",
		"10010111",
		"10011001",
		"10011010",
		"10011001",
		"10011011",
		"10010011",
		"00100001",
		"00001100",
		"00010110",
		"00010100",
		"00100111",
		"00110011",
		"00111101",
		"01000010",
		"01000010",
		"01000110",
		"01001001",
		"01001101",
		"01010000",
		"01010010",
		"01010001",
		"01010010",
		"01010100",
		"01010111",
		"01011010",
		"01011100",
		"01100000",
		"01100010",
		"01100111",
		"01100111",
		"01100010",
		"01011010",
		"01010010",
		"01001100",
		"01000001",
		"00011110",
		"00100011",
		"00101011",
		"00101110",
		"00110001",
		"00101101",
		"00101011",
		"00100011",
		"00011011",
		"00100001",
		"00101010",
		"00011110",
		"00100110",
		"00110000",
		"00110011",
		"01010010",
		"01001010",
		"01010101",
		"01100011",
		"01000001",
		"00101101",
		"01001001",
		"01100111",
		"10010000",
		"10001110",
		"10011001",
		"10101001",
		"10100111",
		"10100110",
		"10100110",
		"10100111",
		"10101011",
		"10101111",
		"10101111",
		"10110001",
		"10110010",
		"10110010",
		"10101111",
		"10100111",
		"10100001",
		"10100010",
		"10100100",
		"10100100",
		"10100011",
		"10011101",
		"10010101",
		"10010001",
		"10001100",
		"10000001",
		"01001011",
		"00011010",
		"00010001",
		"00010011",
		"00010010",
		"00011100",
		"01000010",
		"01010110",
		"01100011",
		"01101110",
		"01110001",
		"01101111",
		"01101101",
		"01100111",
		"01101001",
		"01110101",
		"01110110",
		"01101110",
		"01100010",
		"01100000",
		"01100101",
		"01101110",
		"01111000",
		"01111100",
		"01111010",
		"01110010",
		"01110100",
		"01110010",
		"01110100",
		"01111011",
		"01111110",
		"10000110",
		"10001111",
		"10001110",
		"10010000",
		"10010010",
		"10010001",
		"10010010",
		"10001100",
		"10000101",
		"01110111",
		"01101101",
		"01100111",
		"01101010",
		"01101111",
		"01110100",
		"01111011",
		"01111011",
		"01111001",
		"01111110",
		"01111111",
		"10000000",
		"01111110",
		"10000000",
		"10000011",
		"10001001",
		"10001011",
		"10001101",
		"10001110",
		"10001100",
		"10001100",
		"10001011",
		"10010001",
		"10010101",
		"10010011",
		"10010001",
		"10010111",
		"10010111",
		"10011000",
		"10011011",
		"10100000",
		"10000110",
		"00010110",
		"00001100",
		"00010110",
		"00010010",
		"00011110",
		"00110100",
		"00111100",
		"01000100",
		"01000011",
		"01000011",
		"01000111",
		"01001110",
		"01010010",
		"01010011",
		"01010010",
		"01010011",
		"01010001",
		"01010011",
		"01010110",
		"01011001",
		"01011011",
		"01011101",
		"01011110",
		"01100000",
		"01100000",
		"01011001",
		"01010001",
		"01001010",
		"00111111",
		"00010101",
		"00010101",
		"00010011",
		"00010111",
		"00010111",
		"00010111",
		"00011011",
		"00011101",
		"00011110",
		"00100111",
		"00110010",
		"00100110",
		"00101001",
		"00110111",
		"00110101",
		"00111010",
		"01000110",
		"01001010",
		"00110110",
		"00101010",
		"00011011",
		"00001111",
		"01011101",
		"10010111",
		"10010001",
		"10011100",
		"10101000",
		"10100111",
		"10100110",
		"10100110",
		"10100111",
		"10101011",
		"10101110",
		"10110000",
		"10110001",
		"10110011",
		"10110010",
		"10101110",
		"10101000",
		"10100001",
		"10100001",
		"10100100",
		"10100010",
		"10100001",
		"10011100",
		"10010111",
		"10010100",
		"10001110",
		"01111011",
		"00111100",
		"00011000",
		"00010001",
		"00010010",
		"00010100",
		"00010011",
		"00101101",
		"01001000",
		"01010000",
		"01011100",
		"01101100",
		"01110010",
		"01110100",
		"01101111",
		"01101011",
		"01110011",
		"01110111",
		"01110000",
		"01100010",
		"01011101",
		"01100100",
		"01110010",
		"01111010",
		"01111111",
		"01111011",
		"01110101",
		"01110001",
		"01101010",
		"01101111",
		"01110001",
		"01110111",
		"10000001",
		"10001010",
		"10001001",
		"10001100",
		"10001101",
		"10001111",
		"10010000",
		"10001011",
		"10000101",
		"01110010",
		"01100110",
		"01100011",
		"01101001",
		"01101011",
		"01110000",
		"01111001",
		"01111110",
		"01111011",
		"10000001",
		"10000010",
		"10000001",
		"10000000",
		"10000001",
		"10000101",
		"10000110",
		"10000111",
		"10000100",
		"10001001",
		"10001011",
		"10001100",
		"10001001",
		"10001101",
		"10010010",
		"10010001",
		"10010100",
		"10011001",
		"10011001",
		"10011011",
		"10011110",
		"10100011",
		"01110100",
		"00001101",
		"00001010",
		"00010000",
		"00010100",
		"00010011",
		"00110001",
		"00111101",
		"01000001",
		"01000101",
		"01000111",
		"01000110",
		"01001010",
		"01001111",
		"01010001",
		"01010100",
		"01010011",
		"01010011",
		"01010011",
		"01010111",
		"01011000",
		"01011001",
		"01010111",
		"01011000",
		"01011010",
		"01011010",
		"01010100",
		"01001101",
		"01000111",
		"00111110",
		"00011001",
		"00010100",
		"00001111",
		"00001101",
		"00001100",
		"00001001",
		"00010101",
		"00100100",
		"00101100",
		"00110011",
		"00110111",
		"00111000",
		"00110010",
		"00101000",
		"00111000",
		"01000011",
		"00111010",
		"00101000",
		"00100101",
		"00101001",
		"00011101",
		"00011100",
		"01111000",
		"10010111",
		"10010010",
		"10011011",
		"10100111",
		"10101000",
		"10100101",
		"10100111",
		"10100111",
		"10101100",
		"10101111",
		"10110000",
		"10110010",
		"10110010",
		"10110001",
		"10110000",
		"10101001",
		"10011111",
		"10100010",
		"10100110",
		"10100110",
		"10100100",
		"10011101",
		"10011001",
		"10010100",
		"10010000",
		"01110101",
		"00110010",
		"00010011",
		"00010011",
		"00010011",
		"00010011",
		"00010011",
		"00011001",
		"00111010",
		"01001001",
		"01001101",
		"01011000",
		"01101001",
		"01110100",
		"01110110",
		"01110001",
		"01110000",
		"01110111",
		"01110101",
		"01101100",
		"01100000",
		"01100010",
		"01101111",
		"01111000",
		"01111010",
		"01111001",
		"01110111",
		"01110000",
		"01101001",
		"01101000",
		"01101110",
		"01110011",
		"01111011",
		"10001011",
		"10001100",
		"10001100",
		"10001111",
		"10010010",
		"10001101",
		"10001000",
		"10000000",
		"01110010",
		"01100010",
		"01100010",
		"01100101",
		"01101011",
		"01101100",
		"01110000",
		"01111000",
		"01111000",
		"01111010",
		"01111100",
		"01111110",
		"01111100",
		"01111110",
		"10000100",
		"10000101",
		"10000011",
		"10000011",
		"10000111",
		"10001101",
		"10001100",
		"10001010",
		"10001101",
		"10010011",
		"10010010",
		"10010110",
		"10011001",
		"10011100",
		"10100010",
		"10100001",
		"10100010",
		"01101110",
		"00001010",
		"00001011",
		"00001101",
		"00010101",
		"00001110",
		"00011100",
		"00111011",
		"00111110",
		"01000100",
		"01000111",
		"01001001",
		"01001000",
		"01001010",
		"01001100",
		"01010000",
		"01010001",
		"01010011",
		"01010100",
		"01010101",
		"01010111",
		"01010110",
		"01010011",
		"01010110",
		"01010101",
		"01010100",
		"01010000",
		"01001010",
		"01000100",
		"00111111",
		"00100110",
		"00100110",
		"00100010",
		"00011101",
		"00010100",
		"00001101",
		"00001010",
		"00010111",
		"00100100",
		"00101000",
		"00101001",
		"00101101",
		"00101111",
		"00110010",
		"01010111",
		"01001111",
		"00101111",
		"00011100",
		"00110110",
		"00110110",
		"00101011",
		"00101010",
		"10001011",
		"10010111",
		"10010011",
		"10011010",
		"10100111",
		"10101010",
		"10100101",
		"10100110",
		"10101010",
		"10101101",
		"10101111",
		"10110000",
		"10110001",
		"10110000",
		"10110010",
		"10101111",
		"10100111",
		"10100000",
		"10100100",
		"10100111",
		"10101010",
		"10101000",
		"10100000",
		"10011011",
		"10010101",
		"10010000",
		"01100111",
		"00100110",
		"00010000",
		"00010001",
		"00010010",
		"00010001",
		"00010011",
		"00010011",
		"00100001",
		"01000010",
		"01001010",
		"01001100",
		"01011000",
		"01100111",
		"01110101",
		"01110011",
		"01101010",
		"01101111",
		"01111001",
		"01110111",
		"01101000",
		"01100000",
		"01100111",
		"01110110",
		"01111100",
		"01111100",
		"01111011",
		"01111010",
		"01110000",
		"01101100",
		"01101101",
		"01110000",
		"01110111",
		"01111101",
		"10000111",
		"10001010",
		"10001011",
		"10001011",
		"10001010",
		"10000100",
		"01111000",
		"01101000",
		"01011110",
		"01011101",
		"01100100",
		"01100110",
		"01100100",
		"01101011",
		"01101111",
		"01101110",
		"01101110",
		"01110011",
		"01111000",
		"01110111",
		"01111101",
		"10000001",
		"10000010",
		"10000100",
		"10001001",
		"10001001",
		"10001101",
		"10001100",
		"10001101",
		"10010001",
		"10011000",
		"10010110",
		"10011000",
		"10011100",
		"10011101",
		"10100001",
		"10100100",
		"10100100",
		"01101100",
		"00001001",
		"00001101",
		"00001111",
		"00010101",
		"00011010",
		"00001011",
		"00100000",
		"00111011",
		"01000110",
		"01000111",
		"01001010",
		"01001011",
		"01001100",
		"01001110",
		"01010000",
		"01010001",
		"01010010",
		"01010101",
		"01010011",
		"01010011",
		"01010101",
		"01010011",
		"01010011",
		"01010001",
		"01010000",
		"01001100",
		"01000101",
		"00111110",
		"00111010",
		"00110010",
		"00111100",
		"01000000",
		"01000010",
		"00111010",
		"00101100",
		"00011100",
		"00001111",
		"00010100",
		"00011100",
		"00011110",
		"00100010",
		"00100100",
		"00100101",
		"00100101",
		"00010101",
		"00010110",
		"00110111",
		"01010100",
		"01001100",
		"00101101",
		"00111101",
		"10010110",
		"10010111",
		"10010000",
		"10011011",
		"10100101",
		"10101001",
		"10100110",
		"10100111",
		"10101011",
		"10101101",
		"10101111",
		"10110001",
		"10110001",
		"10110001",
		"10110000",
		"10101101",
		"10100101",
		"10100001",
		"10100100",
		"10101011",
		"10101101",
		"10101010",
		"10100010",
		"10011011",
		"10010111",
		"10010000",
		"01010101",
		"00011100",
		"00010000",
		"00010010",
		"00010010",
		"00010100",
		"00010100",
		"00010001",
		"00011001",
		"00110110",
		"01000110",
		"01001100",
		"01010001",
		"01011100",
		"01101010",
		"01101101",
		"01100110",
		"01100010",
		"01101101",
		"01110011",
		"01110001",
		"01100001",
		"01100000",
		"01101100",
		"01111001",
		"01111101",
		"01111100",
		"01111110",
		"01111011",
		"01110101",
		"01101000",
		"01101000",
		"01101110",
		"01110111",
		"01111011",
		"10000011",
		"10001001",
		"10000111",
		"10001100",
		"10000110",
		"01111001",
		"01100111",
		"01011101",
		"01011110",
		"01100011",
		"01100011",
		"01100110",
		"01101110",
		"01110100",
		"01110011",
		"01101100",
		"01101100",
		"01110011",
		"01110101",
		"01111010",
		"01111110",
		"10000001",
		"10000101",
		"10000100",
		"10001001",
		"10010001",
		"10001110",
		"10001111",
		"10010011",
		"10011000",
		"10011011",
		"10011001",
		"10011011",
		"10011101",
		"10011111",
		"10100010",
		"10100010",
		"01110101",
		"00001110",
		"00001101",
		"00010000",
		"00010110",
		"00100001",
		"00010000",
		"00001011",
		"00011011",
		"00111010",
		"01001001",
		"01001011",
		"01001101",
		"01001110",
		"01001111",
		"01001110",
		"01001110",
		"01001110",
		"01001101",
		"01001110",
		"01010001",
		"01010000",
		"01001110",
		"01001101",
		"01001011",
		"01000111",
		"01000010",
		"00111111",
		"00111011",
		"00111000",
		"00101111",
		"01000110",
		"01001101",
		"01001111",
		"01010111",
		"01001110",
		"01000000",
		"00110010",
		"00100001",
		"00010100",
		"00010100",
		"00011000",
		"00011100",
		"00011101",
		"00011001",
		"00010101",
		"00010111",
		"00011111",
		"00100001",
		"00100111",
		"00011000",
		"01010011",
		"10011011",
		"10011000",
		"10010000",
		"10011100",
		"10100001",
		"10100101",
		"10100011",
		"10100111",
		"10101011",
		"10101101",
		"10110000",
		"10110001",
		"10110001",
		"10110001",
		"10101111",
		"10101001",
		"10100011",
		"10101000",
		"10101110",
		"10101101",
		"10101101",
		"10101011",
		"10100101",
		"10011110",
		"10011010",
		"10001011",
		"01000000",
		"00010010",
		"00010001",
		"00010011",
		"00010010",
		"00010011",
		"00010011",
		"00010011",
		"00010100",
		"00100110",
		"00111101",
		"01001000",
		"01010101",
		"01011001",
		"01100110",
		"01110001",
		"01101000",
		"01100010",
		"01100101",
		"01101101",
		"01110101",
		"01101110",
		"01011110",
		"01011110",
		"01101100",
		"01110111",
		"01111101",
		"01111100",
		"01111111",
		"01110101",
		"01101111",
		"01101100",
		"01101011",
		"01110001",
		"01111001",
		"01111111",
		"10000010",
		"10001000",
		"10001110",
		"10001110",
		"10000101",
		"01110010",
		"01100111",
		"01100001",
		"01100001",
		"01100001",
		"01101010",
		"01110100",
		"01111001",
		"01110110",
		"01110011",
		"01110100",
		"01111000",
		"01110100",
		"01110011",
		"01110110",
		"01111011",
		"01111110",
		"10000001",
		"10001010",
		"10001111",
		"10001101",
		"10001111",
		"10010011",
		"10011010",
		"10011010",
		"10011010",
		"10011010",
		"10011101",
		"10011101",
		"10011110",
		"10100000",
		"01111001",
		"00010001",
		"00001101",
		"00010010",
		"00011011",
		"00100111",
		"00100011",
		"00010100",
		"00001101",
		"00010010",
		"00101010",
		"00111111",
		"01001101",
		"01010011",
		"01010001",
		"01010000",
		"01001110",
		"01010000",
		"01001101",
		"01001100",
		"01001100",
		"01001010",
		"01000111",
		"01000001",
		"01000000",
		"00111110",
		"00111110",
		"00111111",
		"00111101",
		"00111010",
		"00101101",
		"01000100",
		"01001001",
		"01010111",
		"01101000",
		"01100011",
		"01010101",
		"01001001",
		"01000111",
		"00111011",
		"00100111",
		"00010111",
		"00010011",
		"00010011",
		"00010011",
		"00010100",
		"00011110",
		"00100100",
		"00100011",
		"00100001",
		"00100001",
		"01110010",
		"10011110",
		"10011001",
		"10001110",
		"10011101",
		"10100000",
		"10100000",
		"10100001",
		"10101000",
		"10101101",
		"10101101",
		"10110000",
		"10110010",
		"10110011",
		"10110101",
		"10110111",
		"10110011",
		"10101000",
		"10101110",
		"10110011",
		"10110001",
		"10101111",
		"10101011",
		"10100011",
		"10011110",
		"10011101",
		"01111110",
		"00101011",
		"00001111",
		"00010011",
		"00010001",
		"00010001",
		"00010010",
		"00010010",
		"00010011",
		"00010100",
		"00011101",
		"00110100",
		"01000001",
		"01001111",
		"01011011",
		"01100011",
		"01101101",
		"01101101",
		"01100110",
		"01100110",
		"01101111",
		"01110100",
		"01110001",
		"01101000",
		"01011100",
		"01011111",
		"01101010",
		"01110110",
		"01111011",
		"01111110",
		"01111001",
		"01110010",
		"01101100",
		"01100100",
		"01101010",
		"01110100",
		"01111100",
		"10000100",
		"10001010",
		"10001100",
		"10001110",
		"10000110",
		"01110110",
		"01100111",
		"01100100",
		"01011110",
		"01100000",
		"01101001",
		"01110011",
		"01111000",
		"01111000",
		"01111101",
		"10000011",
		"10000010",
		"10000010",
		"01111101",
		"01111101",
		"01111110",
		"10000011",
		"10000110",
		"10001000",
		"10001001",
		"10001101",
		"10010010",
		"10010010",
		"10010111",
		"10011011",
		"10011000",
		"10011011",
		"10011101",
		"10011100",
		"10011101",
		"10011111",
		"01110001",
		"00001100",
		"00001101",
		"00010100",
		"00100101",
		"00111110",
		"00111100",
		"00101100",
		"00011100",
		"00001110",
		"00001100",
		"00010000",
		"00011110",
		"00110001",
		"00111111",
		"01000101",
		"01000110",
		"01000111",
		"01000111",
		"01000100",
		"01000001",
		"00111101",
		"00111011",
		"00111010",
		"00111101",
		"00111110",
		"01000100",
		"01000100",
		"00111110",
		"00111010",
		"00111010",
		"01001100",
		"01000110",
		"01001001",
		"01001101",
		"01001110",
		"01001100",
		"01000100",
		"01000000",
		"01000001",
		"01000000",
		"00110010",
		"00011011",
		"00001101",
		"00001100",
		"00010000",
		"00010110",
		"00011010",
		"00011101",
		"00011001",
		"00100001",
		"10000110",
		"10011111",
		"10011101",
		"10001111",
		"10011110",
		"10100000",
		"10100001",
		"10100010",
		"10100111",
		"10101100",
		"10101110",
		"10101111",
		"10110010",
		"10110001",
		"10110100",
		"10110011",
		"10101110",
		"10101001",
		"10110001",
		"10110011",
		"10110001",
		"10101111",
		"10101100",
		"10100100",
		"10011111",
		"10011101",
		"01100010",
		"00010111",
		"00001111",
		"00010011",
		"00010001",
		"00010010",
		"00010010",
		"00010011",
		"00010100",
		"00010100",
		"00011000",
		"00101010",
		"00111110",
		"01000110",
		"01011011",
		"01100010",
		"01100111",
		"01100110",
		"01101010",
		"01101011",
		"01101111",
		"01110100",
		"01110100",
		"01101000",
		"01010110",
		"01010110",
		"01100001",
		"01101110",
		"01110111",
		"01110111",
		"01110111",
		"01110011",
		"01101001",
		"01100100",
		"01101001",
		"01101101",
		"01110111",
		"10000000",
		"10000111",
		"10001001",
		"10001001",
		"10001000",
		"01110001",
		"01100001",
		"01100100",
		"01100110",
		"01100100",
		"01100111",
		"01110001",
		"01110011",
		"01110101",
		"01111100",
		"10000100",
		"10000101",
		"10000100",
		"10000101",
		"10001000",
		"10000100",
		"10000110",
		"10001001",
		"10001010",
		"10001101",
		"10001101",
		"10010010",
		"10010001",
		"10010101",
		"10011011",
		"10011111",
		"10011110",
		"10011001",
		"10011100",
		"10011110",
		"10100000",
		"01100101",
		"00000111",
		"00001101",
		"00010011",
		"00100101",
		"01000100",
		"01010011",
		"01001001",
		"00111001",
		"00010100",
		"00001100",
		"00001010",
		"00001001",
		"00001010",
		"00010000",
		"00011000",
		"00100011",
		"00101111",
		"00110110",
		"00110110",
		"00111100",
		"00111101",
		"00111101",
		"00111101",
		"00111100",
		"00111110",
		"00111111",
		"00111111",
		"01000001",
		"00111101",
		"01010000",
		"01101101",
		"01100011",
		"01011011",
		"01011000",
		"01010001",
		"01001110",
		"01000111",
		"00111011",
		"00110100",
		"00110100",
		"00101110",
		"00100011",
		"00010111",
		"00001101",
		"00001110",
		"00010011",
		"00011000",
		"00011001",
		"00010011",
		"00110100",
		"10011000",
		"10011101",
		"10011011",
		"10001110",
		"10011110",
		"10100010",
		"10100011",
		"10100110",
		"10101000",
		"10101011",
		"10101101",
		"10101111",
		"10110000",
		"10110001",
		"10110000",
		"10101100",
		"10100101",
		"10100101",
		"10101100",
		"10110001",
		"10110001",
		"10110001",
		"10101110",
		"10100111",
		"10100010",
		"10010010",
		"00111010",
		"00001110",
		"00010001",
		"00010010",
		"00010011",
		"00010011",
		"00010011",
		"00010100",
		"00010100",
		"00010110",
		"00010100",
		"00100100",
		"00111111",
		"01000101",
		"01010010",
		"01100000",
		"01101010",
		"01100111",
		"01100101",
		"01101101",
		"01101110",
		"01110011",
		"01110110",
		"01101000",
		"01010111",
		"01010101",
		"01011101",
		"01101000",
		"01110011",
		"01110110",
		"01111000",
		"01111000",
		"01101100",
		"01100111",
		"01100010",
		"01100100",
		"01110000",
		"01111100",
		"10000100",
		"10000010",
		"10000000",
		"01111000",
		"01100110",
		"01011011",
		"01011011",
		"01100011",
		"01101001",
		"01100110",
		"01101111",
		"01110000",
		"01110100",
		"01111100",
		"10000000",
		"10000010",
		"10000100",
		"10000110",
		"10001010",
		"10001010",
		"10001010",
		"10001110",
		"10010000",
		"10010010",
		"10001111",
		"10010011",
		"10010011",
		"10010111",
		"10011111",
		"10100010",
		"10011110",
		"10011010",
		"10011111",
		"10011101",
		"10011111",
		"01001111",
		"00000101",
		"00001011",
		"00001101",
		"00010110",
		"00101111",
		"01001100",
		"01010000",
		"01111011",
		"01000001",
		"00001001",
		"00001011",
		"00001011",
		"00010001",
		"00011101",
		"00100110",
		"00110001",
		"00111011",
		"00111100",
		"00111100",
		"01000000",
		"01000000",
		"01000010",
		"01000000",
		"00111110",
		"00111111",
		"00111101",
		"00111110",
		"01000010",
		"00111110",
		"01001111",
		"01101110",
		"01100100",
		"01100011",
		"01100001",
		"01011111",
		"01011011",
		"01011010",
		"01010101",
		"01010001",
		"01010000",
		"01001011",
		"01001110",
		"01001100",
		"01001001",
		"01000110",
		"01001001",
		"01001000",
		"01000100",
		"00110111",
		"01100011",
		"10011101",
		"10011111",
		"10011000",
		"10001110",
		"10011110",
		"10100011",
		"10100001",
		"10100101",
		"10101001",
		"10101010",
		"10101011",
		"10101110",
		"10101111",
		"10110000",
		"10110001",
		"10101101",
		"10101000",
		"10101000",
		"10101110",
		"10110010",
		"10110011",
		"10101111",
		"10101101",
		"10101000",
		"10100011",
		"01101110",
		"00011011",
		"00001110",
		"00010001",
		"00010001",
		"00010011",
		"00010010",
		"00010101",
		"00010110",
		"00010111",
		"00010110",
		"00011000",
		"00100100",
		"01000000",
		"01000110",
		"01001111",
		"01011001",
		"01100100",
		"01100110",
		"01100000",
		"01101000",
		"01110010",
		"01110100",
		"01101101",
		"01011111",
		"01010110",
		"01010100",
		"01010111",
		"01100010",
		"01101010",
		"01110111",
		"01111001",
		"01110111",
		"01101111",
		"01101000",
		"01100110",
		"01100101",
		"01110000",
		"01111001",
		"10000000",
		"01111101",
		"01111001",
		"01110011",
		"01100001",
		"01010111",
		"01010110",
		"01011110",
		"01100100",
		"01101011",
		"01101110",
		"01110010",
		"01110111",
		"01111111",
		"10000001",
		"10000010",
		"10000110",
		"10001010",
		"10001011",
		"10001110",
		"10001101",
		"10010000",
		"10010001",
		"10010011",
		"10010001",
		"10010010",
		"10010010",
		"10011001",
		"10100001",
		"10100000",
		"10011100",
		"10011001",
		"10011011",
		"10011011",
		"10011001",
		"00110010",
		"00000101",
		"00001010",
		"00001100",
		"00001100",
		"00010101",
		"00100101",
		"00110001",
		"01010101",
		"01110111",
		"00010000",
		"00001011",
		"00001111",
		"00011100",
		"00101010",
		"00110000",
		"00110111",
		"00111101",
		"01000001",
		"01000011",
		"01000011",
		"01000100",
		"01000010",
		"01000000",
		"00111111",
		"01000000",
		"00111110",
		"00111100",
		"00111101",
		"00111010",
		"01101001",
		"10010101",
		"10001101",
		"10001010",
		"10000100",
		"01111011",
		"01110100",
		"01101101",
		"01100111",
		"01100010",
		"01011110",
		"01011010",
		"01011100",
		"01011011",
		"01010111",
		"01010011",
		"01010011",
		"01010000",
		"01001001",
		"01000110",
		"01111111",
		"10011111",
		"10011110",
		"10001101",
		"10010001",
		"10011101",
		"10100000",
		"10100010",
		"10100010",
		"10100110",
		"10101011",
		"10101101",
		"10101110",
		"10101111",
		"10101111",
		"10101111",
		"10101100",
		"10101010",
		"10101101",
		"10110001",
		"10110100",
		"10110010",
		"10110000",
		"10101101",
		"10100110",
		"10010110",
		"00111110",
		"00001110",
		"00010000",
		"00010000",
		"00010001",
		"00010011",
		"00010010",
		"00010100",
		"00010110",
		"00010111",
		"00011000",
		"00011000",
		"00011100",
		"00110100",
		"01000000",
		"01001010",
		"01010100",
		"01011000",
		"01011011",
		"01011001",
		"01011110",
		"01101001",
		"01110010",
		"01101001",
		"01011000",
		"01010011",
		"01100000",
		"01011100",
		"01100010",
		"01101111",
		"01111000",
		"01111010",
		"01110011",
		"01101101",
		"01100101",
		"01100101",
		"01101001",
		"01110001",
		"01110110",
		"01111100",
		"01111100",
		"01111010",
		"01110010",
		"01011100",
		"01010010",
		"01010110",
		"01011001",
		"01011101",
		"01101010",
		"01101110",
		"01101111",
		"01110111",
		"01111101",
		"01111110",
		"10000011",
		"10000101",
		"10001000",
		"10000111",
		"10001011",
		"10001010",
		"10001000",
		"10001111",
		"10010001",
		"10010010",
		"10010010",
		"10010010",
		"10010111",
		"10011100",
		"10011100",
		"10011011",
		"10011001",
		"10010111",
		"10011001",
		"10001000",
		"00010111",
		"00001000",
		"00001010",
		"00001010",
		"00001010",
		"00001011",
		"00001110",
		"00010010",
		"00010000",
		"00100111",
		"00010100",
		"00001001",
		"00010011",
		"00100010",
		"00101110",
		"00110111",
		"00111100",
		"01000000",
		"01000110",
		"01001010",
		"01001010",
		"01000111",
		"01000101",
		"01000011",
		"01000010",
		"00111110",
		"00111100",
		"00111100",
		"00111101",
		"00111100",
		"01111000",
		"10101110",
		"10100110",
		"10100011",
		"10011101",
		"10010101",
		"10001111",
		"10001000",
		"10000001",
		"01110111",
		"01101110",
		"01101010",
		"01100001",
		"01011110",
		"01011000",
		"01010111",
		"01010110",
		"01010101",
		"01001100",
		"01010101",
		"10001111",
		"10011101",
		"10011010",
		"10000111",
		"10010110",
		"10011011",
		"10011110",
		"10100010",
		"10100100",
		"10101001",
		"10101100",
		"10101111",
		"10110000",
		"10110000",
		"10110000",
		"10101111",
		"10101100",
		"10101011",
		"10101111",
		"10110011",
		"10110100",
		"10110011",
		"10110010",
		"10101110",
		"10101000",
		"01110110",
		"00011100",
		"00001110",
		"00010001",
		"00010001",
		"00010010",
		"00010011",
		"00010101",
		"00010111",
		"00011001",
		"00011010",
		"00011101",
		"00011100",
		"00011101",
		"00100110",
		"00111011",
		"01000001",
		"01010000",
		"01010011",
		"01010111",
		"01011010",
		"01100001",
		"01101000",
		"01110010",
		"01110011",
		"01100011",
		"01011011",
		"01100011",
		"01101000",
		"01101100",
		"01110101",
		"01111011",
		"01111011",
		"01110110",
		"01110000",
		"01101010",
		"01101000",
		"01101100",
		"01110010",
		"01110110",
		"01111110",
		"01111101",
		"01110111",
		"01100111",
		"01011101",
		"01010110",
		"01011101",
		"01011011",
		"01011100",
		"01100010",
		"01101000",
		"01101000",
		"01110011",
		"01111001",
		"01111001",
		"10000000",
		"10000000",
		"10000011",
		"10000110",
		"10001010",
		"10001011",
		"10001000",
		"10001101",
		"10010000",
		"10001101",
		"10001101",
		"10010000",
		"10010110",
		"10011101",
		"10011010",
		"10011011",
		"10011001",
		"10010111",
		"10011010",
		"01011001",
		"00000101",
		"00001011",
		"00001011",
		"00001011",
		"00001011",
		"00001100",
		"00001011",
		"00001100",
		"00001100",
		"00001100",
		"00001101",
		"00001011",
		"00010101",
		"00101010",
		"00110101",
		"00111010",
		"01000100",
		"01001011",
		"01001101",
		"01001010",
		"01001000",
		"01000111",
		"01000100",
		"01000011",
		"01000000",
		"00111101",
		"00111011",
		"00111101",
		"01000000",
		"00111111",
		"01111111",
		"10111001",
		"10110001",
		"10101111",
		"10101011",
		"10100101",
		"10011111",
		"10011001",
		"10010100",
		"10001011",
		"10000010",
		"01111011",
		"01110010",
		"01100111",
		"01011110",
		"01010111",
		"01010011",
		"01010000",
		"01001001",
		"01100111",
		"10010010",
		"10011001",
		"10001101",
		"10001001",
		"10011101",
		"10011100",
		"10011100",
		"10011110",
		"10100101",
		"10101010",
		"10101110",
		"10110001",
		"10110000",
		"10110001",
		"10110001",
		"10101110",
		"10101110",
		"10110000",
		"10110100",
		"10110101",
		"10110110",
		"10110101",
		"10110101",
		"10101111",
		"10100010",
		"01000101",
		"00001011",
		"00001111",
		"00010011",
		"00010100",
		"00010011",
		"00010101",
		"00010111",
		"00011000",
		"00011001",
		"00011110",
		"00011111",
		"00011111",
		"00011110",
		"00100001",
		"00110100",
		"00111110",
		"01001111",
		"01011001",
		"01011010",
		"01010110",
		"01011100",
		"01100111",
		"01110001",
		"01110001",
		"01100111",
		"01011100",
		"01011101",
		"01101001",
		"01101100",
		"01110011",
		"01111010",
		"01111111",
		"01111000",
		"01110000",
		"01101110",
		"01101110",
		"01110001",
		"01110110",
		"01111101",
		"01111111",
		"01111011",
		"01110000",
		"01100010",
		"01011100",
		"01010101",
		"01011110",
		"01011100",
		"01010111",
		"01011101",
		"01011111",
		"01100100",
		"01101001",
		"01100111",
		"01101110",
		"01110100",
		"01111001",
		"10000000",
		"10000100",
		"10001000",
		"10001001",
		"10001000",
		"10001011",
		"10001110",
		"10001010",
		"10001011",
		"10001111",
		"10011001",
		"10100000",
		"10011100",
		"10011011",
		"10010111",
		"10010011",
		"10001100",
		"00101001",
		"00000111",
		"00001011",
		"00001100",
		"00001010",
		"00001010",
		"00001011",
		"00001100",
		"00001011",
		"00001011",
		"00001100",
		"00001100",
		"00001100",
		"00010100",
		"00101001",
		"00110110",
		"00111101",
		"01000110",
		"01010000",
		"01001101",
		"01001100",
		"01001001",
		"01000101",
		"01000010",
		"01000000",
		"00111110",
		"00111011",
		"00111100",
		"00111110",
		"01000100",
		"01000101",
		"10000110",
		"10111100",
		"10110110",
		"10110100",
		"10110001",
		"10101101",
		"10100110",
		"10100001",
		"10011101",
		"10010111",
		"10010000",
		"10001101",
		"10000011",
		"01110000",
		"01100100",
		"01010111",
		"01001111",
		"01001010",
		"01000101",
		"01111011",
		"10010000",
		"10010101",
		"10000110",
		"10001100",
		"10011011",
		"10011001",
		"10011010",
		"10011110",
		"10100100",
		"10101011",
		"10101111",
		"10110000",
		"10110000",
		"10110010",
		"10110000",
		"10101101",
		"10101111",
		"10110011",
		"10110110",
		"10110111",
		"10110111",
		"10110101",
		"10110010",
		"10101110",
		"10001100",
		"00011100",
		"00001111",
		"00010011",
		"00010101",
		"00010110",
		"00011000",
		"00011001",
		"00011001",
		"00011101",
		"00011101",
		"00011110",
		"00011110",
		"00011111",
		"00100011",
		"00100100",
		"00101010",
		"00111001",
		"01000100",
		"01010011",
		"01011010",
		"01010110",
		"01011100",
		"01100100",
		"01101101",
		"01110011",
		"01100110",
		"01011011",
		"01011110",
		"01101001",
		"01110000",
		"01110011",
		"01111010",
		"10000000",
		"01111101",
		"01110111",
		"01110100",
		"01110010",
		"01110011",
		"01110111",
		"01111100",
		"01111111",
		"01111010",
		"01101110",
		"01100011",
		"01010000",
		"01001010",
		"01010011",
		"01010100",
		"01001100",
		"01001101",
		"01001101",
		"01010100",
		"01010111",
		"01011000",
		"01011110",
		"01100111",
		"01110001",
		"01111010",
		"10000001",
		"10000101",
		"10000101",
		"10001001",
		"10001010",
		"10001100",
		"10001011",
		"10001110",
		"10010101",
		"10011111",
		"10011101",
		"10011001",
		"10010111",
		"10010110",
		"10000110",
		"00111111",
		"00000101",
		"00001000",
		"00001010",
		"00001100",
		"00001001",
		"00000110",
		"00000101",
		"00000100",
		"00000111",
		"00001001",
		"00001010",
		"00001011",
		"00001010",
		"00001110",
		"00100101",
		"00110100",
		"00111011",
		"01000011",
		"01000101",
		"01000111",
		"01001000",
		"01001000",
		"01000011",
		"01000001",
		"01000000",
		"00111110",
		"01000000",
		"01000001",
		"01000110",
		"01001001",
		"01000101",
		"10001001",
		"10111101",
		"10110111",
		"10110101",
		"10110101",
		"10110011",
		"10101101",
		"10100111",
		"10100100",
		"10011101",
		"10010111",
		"10010000",
		"10001001",
		"01111001",
		"01101111",
		"01011111",
		"01010100",
		"01001000",
		"01010100",
		"10000111",
		"10010000",
		"10001101",
		"10000100",
		"10010100",
		"10011010",
		"10010111",
		"10011010",
		"10011110",
		"10100100",
		"10101101",
		"10110000",
		"10110001",
		"10110010",
		"10110010",
		"10110000",
		"10110000",
		"10110010",
		"10110101",
		"10110111",
		"10111000",
		"10110111",
		"10110101",
		"10110010",
		"10101111",
		"01011010",
		"00001111",
		"00010101",
		"00010111",
		"00011001",
		"00011011",
		"00011011",
		"00011010",
		"00011100",
		"00011111",
		"00011111",
		"00011110",
		"00100001",
		"00100011",
		"00100000",
		"00100010",
		"00100011",
		"00101111",
		"00111100",
		"01000110",
		"01001111",
		"01010000",
		"01011010",
		"01100011",
		"01101010",
		"01110100",
		"01101111",
		"01011001",
		"01011000",
		"01100100",
		"01101010",
		"01110110",
		"01111100",
		"10000001",
		"10000001",
		"01111011",
		"01110110",
		"01110010",
		"01110010",
		"01110101",
		"01111000",
		"01111100",
		"01111011",
		"01110101",
		"01101110",
		"01010101",
		"01000101",
		"01000110",
		"01001010",
		"01001001",
		"01000110",
		"01001011",
		"01001100",
		"01010001",
		"01010110",
		"01011001",
		"01100101",
		"01110001",
		"01110101",
		"01111010",
		"01111111",
		"10000001",
		"10000100",
		"10001001",
		"10001011",
		"10001010",
		"10001110",
		"10010111",
		"10011010",
		"10011001",
		"10011001",
		"10010110",
		"10001010",
		"01001111",
		"00100011",
		"00101110",
		"01000110",
		"01001100",
		"01001011",
		"01001100",
		"01000011",
		"00110011",
		"00100011",
		"00010100",
		"00001000",
		"00000100",
		"00000110",
		"00000111",
		"00001000",
		"00010100",
		"00101011",
		"00110100",
		"00111100",
		"01000001",
		"01000001",
		"01000010",
		"01000010",
		"01000001",
		"01000001",
		"01000011",
		"01000010",
		"01000011",
		"01000111",
		"01001001",
		"01001100",
		"01001001",
		"10001010",
		"11000001",
		"10111010",
		"10111000",
		"10110110",
		"10110101",
		"10110101",
		"10110001",
		"10101000",
		"10100100",
		"10011110",
		"10010110",
		"10001100",
		"10000001",
		"01110010",
		"01100100",
		"01010010",
		"01000110",
		"01100111",
		"10001001",
		"10001100",
		"10000101",
		"10000110",
		"10011010",
		"10011010",
		"10011010",
		"10011100",
		"10011111",
		"10100100",
		"10101100",
		"10110000",
		"10110011",
		"10110011",
		"10110010",
		"10110000",
		"10101111",
		"10110010",
		"10110101",
		"10110111",
		"10110111",
		"10110110",
		"10110101",
		"10110101",
		"10010111",
		"00100010",
		"00010001",
		"00010110",
		"00011000",
		"00011010",
		"00011100",
		"00011101",
		"00011100",
		"00011100",
		"00011111",
		"00011111",
		"00011111",
		"00100001",
		"00100001",
		"00011111",
		"00100010",
		"00100000",
		"00100101",
		"00110101",
		"01000000",
		"01000111",
		"01000111",
		"01010001",
		"01011111",
		"01100111",
		"01110001",
		"01101110",
		"01011110",
		"01010110",
		"01011101",
		"01100110",
		"01101111",
		"01111001",
		"10000110",
		"10000111",
		"10000100",
		"01111010",
		"01110011",
		"01110101",
		"01111001",
		"01111011",
		"01111001",
		"01110111",
		"01110101",
		"01100111",
		"01010110",
		"01000100",
		"01000011",
		"01000100",
		"01000100",
		"01000011",
		"01001001",
		"01001100",
		"01010101",
		"01100001",
		"01100000",
		"01100001",
		"01101010",
		"01110001",
		"01111010",
		"01111110",
		"10000010",
		"10000011",
		"10000101",
		"10001011",
		"10001100",
		"10010001",
		"10010011",
		"10010111",
		"10010110",
		"10010110",
		"10000001",
		"00111110",
		"00100011",
		"01001001",
		"01011010",
		"01100101",
		"01101000",
		"01101000",
		"01101100",
		"01101100",
		"01101000",
		"01100011",
		"01011100",
		"01001001",
		"00110011",
		"00011110",
		"00001101",
		"00000110",
		"00000101",
		"00010010",
		"00100101",
		"00110011",
		"00111010",
		"00111101",
		"00111111",
		"01000000",
		"01000011",
		"01000011",
		"01000110",
		"01000101",
		"01000111",
		"01001101",
		"01001101",
		"01010000",
		"01001011",
		"10010000",
		"11001000",
		"11000100",
		"11001000",
		"11001000",
		"11000101",
		"11000100",
		"10111100",
		"10101111",
		"10100110",
		"10100000",
		"10010111",
		"10001110",
		"10000011",
		"01110001",
		"01011101",
		"01001110",
		"01000110",
		"01110111",
		"10001010",
		"10001000",
		"10000000",
		"10001011",
		"10011010",
		"10010101",
		"10011000",
		"10011011",
		"10011110",
		"10100110",
		"10101100",
		"10101111",
		"10110010",
		"10110011",
		"10110100",
		"10110010",
		"10110000",
		"10110010",
		"10110101",
		"10110110",
		"10110111",
		"10110111",
		"10110111",
		"10110100",
		"01011101",
		"00001110",
		"00010110",
		"00011001",
		"00011010",
		"00011011",
		"00011100",
		"00011110",
		"00011101",
		"00011100",
		"00011111",
		"00011111",
		"00100000",
		"00100000",
		"00011111",
		"00100000",
		"00100001",
		"00011111",
		"00011111",
		"00101010",
		"00111011",
		"01000010",
		"01000100",
		"01001111",
		"01011011",
		"01100010",
		"01101001",
		"01101011",
		"01100000",
		"01010110",
		"01010110",
		"01011111",
		"01100110",
		"01110111",
		"10000001",
		"10000111",
		"10000010",
		"01111001",
		"01110111",
		"01110010",
		"01111001",
		"01111000",
		"01111000",
		"01110111",
		"01110000",
		"01011111",
		"01001111",
		"01000011",
		"01000010",
		"01000000",
		"01000011",
		"01000101",
		"01000111",
		"01001100",
		"01010101",
		"01011100",
		"01011101",
		"01100010",
		"01101110",
		"01111000",
		"10000000",
		"10000111",
		"10000111",
		"10001001",
		"10001011",
		"10001100",
		"10001100",
		"10010000",
		"10010101",
		"10010110",
		"10010011",
		"01110101",
		"00101000",
		"00000110",
		"00101000",
		"01001100",
		"01011011",
		"01101100",
		"01111010",
		"10000100",
		"10001001",
		"10001100",
		"10001010",
		"01111101",
		"01110001",
		"01101011",
		"01100101",
		"01100000",
		"01010101",
		"01000011",
		"00101011",
		"00011000",
		"00010011",
		"00011001",
		"00100011",
		"00110010",
		"00111001",
		"00111110",
		"01000001",
		"01000101",
		"01000111",
		"01001010",
		"01001101",
		"01001111",
		"01010000",
		"01010001",
		"01001100",
		"10011010",
		"11011011",
		"11010111",
		"11010111",
		"11010111",
		"11010101",
		"11001111",
		"10111111",
		"10110011",
		"10101000",
		"10011110",
		"10010101",
		"10000101",
		"01110010",
		"01100010",
		"01010001",
		"00111111",
		"01001001",
		"01111000",
		"10000000",
		"01111111",
		"01111101",
		"10001110",
		"10010011",
		"10010001",
		"10010101",
		"10011001",
		"10011100",
		"10100111",
		"10101110",
		"10110000",
		"10110011",
		"10110100",
		"10110100",
		"10110011",
		"10110010",
		"10110101",
		"10110111",
		"10111010",
		"10111010",
		"10111000",
		"10110111",
		"10010110",
		"00100000",
		"00010001",
		"00010111",
		"00011010",
		"00011010",
		"00011100",
		"00011011",
		"00011101",
		"00011111",
		"00011110",
		"00011110",
		"00100000",
		"00011110",
		"00011100",
		"00100000",
		"00100000",
		"00100001",
		"00100000",
		"00011101",
		"00100011",
		"00110000",
		"00111100",
		"01000011",
		"01001000",
		"01010100",
		"01100001",
		"01101011",
		"01101101",
		"01100101",
		"01011000",
		"01010000",
		"01010100",
		"01011100",
		"01101000",
		"01110010",
		"01111100",
		"01111100",
		"01110111",
		"01110001",
		"01110011",
		"01110011",
		"01110011",
		"01110100",
		"01110010",
		"01011100",
		"01010011",
		"01000101",
		"00111010",
		"00111000",
		"00110100",
		"00111001",
		"00111101",
		"01000010",
		"01000101",
		"01001000",
		"01001110",
		"01010100",
		"01011001",
		"01100111",
		"01110111",
		"01111001",
		"10000000",
		"10001011",
		"10010000",
		"10001100",
		"10001011",
		"10001110",
		"10010011",
		"10010101",
		"10001101",
		"01100100",
		"00011001",
		"00000100",
		"00101011",
		"00110111",
		"01001010",
		"01011011",
		"01101001",
		"10000000",
		"10010110",
		"10100011",
		"10101001",
		"10101010",
		"10011110",
		"10010010",
		"10000011",
		"01110011",
		"01101100",
		"01101101",
		"01101011",
		"01101000",
		"01100000",
		"01010010",
		"01000100",
		"00110001",
		"00100110",
		"00100111",
		"00110010",
		"00111101",
		"01000001",
		"01000111",
		"01001100",
		"01001110",
		"01010000",
		"01010001",
		"01010001",
		"01001010",
		"10011000",
		"11011000",
		"11010100",
		"11010101",
		"11010101",
		"11010110",
		"11010000",
		"10111111",
		"10110000",
		"10100101",
		"10011011",
		"10001101",
		"01110100",
		"01100000",
		"01010000",
		"00111110",
		"00101010",
		"00111101",
		"01100011",
		"01110011",
		"01110000",
		"01110011",
		"10001010",
		"10001011",
		"10001000",
		"10001110",
		"10010100",
		"10011000",
		"10100101",
		"10101110",
		"10110000",
		"10110010",
		"10110100",
		"10110011",
		"10110100",
		"10110100",
		"10110111",
		"10111001",
		"10111001",
		"10111000",
		"10111001",
		"10101111",
		"01000111",
		"00001111",
		"00010101",
		"00011000",
		"00011011",
		"00011101",
		"00011110",
		"00011110",
		"00011110",
		"00100000",
		"00011110",
		"00011110",
		"00011111",
		"00011110",
		"00011110",
		"00011101",
		"00011101",
		"00011101",
		"00011111",
		"00011110",
		"00011101",
		"00100001",
		"00101111",
		"00111101",
		"01000110",
		"01001101",
		"01100000",
		"01101011",
		"01110100",
		"01101001",
		"01010110",
		"01001101",
		"01001100",
		"01010101",
		"01011011",
		"01100101",
		"01101000",
		"01100111",
		"01011111",
		"01100100",
		"01101011",
		"01101110",
		"01101110",
		"01101010",
		"01100111",
		"01011010",
		"01010001",
		"01000110",
		"00111000",
		"00110001",
		"00110010",
		"00110100",
		"00110011",
		"00110110",
		"00111001",
		"00111100",
		"01000100",
		"01000101",
		"01001010",
		"01010000",
		"01100001",
		"01101100",
		"01111000",
		"10000101",
		"10001010",
		"10001010",
		"10000111",
		"10000111",
		"10000001",
		"01101110",
		"00111000",
		"00001000",
		"00001110",
		"01000001",
		"01101101",
		"01001010",
		"01001001",
		"01010110",
		"01101110",
		"10010010",
		"10100101",
		"10101001",
		"10110010",
		"11000011",
		"11000111",
		"11001000",
		"10111110",
		"10100001",
		"10010000",
		"10000111",
		"01111110",
		"01110101",
		"01110111",
		"01110111",
		"01110010",
		"01101101",
		"01100001",
		"01001111",
		"01000110",
		"00111110",
		"00111011",
		"01000000",
		"01000110",
		"01001100",
		"01001100",
		"01001110",
		"01010000",
		"01000111",
		"10010100",
		"11001100",
		"11001000",
		"11000110",
		"11000100",
		"11000010",
		"10111110",
		"10110111",
		"10101011",
		"10011111",
		"10001101",
		"01101111",
		"01010111",
		"01000110",
		"00110100",
		"00100011",
		"00010010",
		"00101000",
		"01001000",
		"01010111",
		"01010101",
		"01010100",
		"01110001",
		"01110100",
		"01110110",
		"01111011",
		"10000101",
		"10010000",
		"10011011",
		"10100111",
		"10101101",
		"10101111",
		"10101110",
		"10101110",
		"10110000",
		"10110011",
		"10110111",
		"10111000",
		"10110111",
		"10110111",
		"10110100",
		"01110000",
		"00010001",
		"00010110",
		"00011000",
		"00011010",
		"00011011",
		"00011100",
		"00011100",
		"00011100",
		"00011100",
		"00011101",
		"00011110",
		"00011110",
		"00011101",
		"00011101",
		"00011100",
		"00011100",
		"00011101",
		"00011100",
		"00011011",
		"00011111",
		"00011101",
		"00011011",
		"00100011",
		"00101111",
		"00111100",
		"01000101",
		"01011010",
		"01101001",
		"01110011",
		"01101100",
		"01011010",
		"01001111",
		"01001101",
		"01001100",
		"01010000",
		"01010100",
		"01010101",
		"01011000",
		"01010111",
		"01011010",
		"01100101",
		"01100100",
		"01100110",
		"01101001",
		"01011111",
		"01010111",
		"01000010",
		"00110101",
		"00100111",
		"00100111",
		"00101010",
		"00101111",
		"00110011",
		"00110011",
		"00110001",
		"00110000",
		"00110011",
		"00111101",
		"00111011",
		"00111010",
		"01000110",
		"01001101",
		"01010101",
		"01011111",
		"01011010",
		"01100010",
		"01110000",
		"10000001",
		"10001110",
		"01111001",
		"01100010",
		"01111011",
		"10001110",
		"01111100",
		"01100100",
		"01100010",
		"01010001",
		"01011110",
		"01110010",
		"10001000",
		"10010011",
		"10011110",
		"10101101",
		"11001001",
		"11010000",
		"11011100",
		"11011101",
		"11011011",
		"11010001",
		"11001000",
		"10111110",
		"10111000",
		"10111000",
		"10111001",
		"10110001",
		"10111001",
		"10100101",
		"10010101",
		"10001000",
		"01100111",
		"01010101",
		"01001010",
		"01000001",
		"01000010",
		"01000101",
		"01001001",
		"01001100",
		"01000110",
		"10001011",
		"11000110",
		"11000000",
		"10111110",
		"10111011",
		"10110111",
		"10110010",
		"10101100",
		"10011111",
		"10010100",
		"10001100",
		"10001000",
		"10001000",
		"10001010",
		"10001101",
		"10001101",
		"10001100",
		"10010100",
		"10011110",
		"10100100",
		"10100110",
		"10100000",
		"10100011",
		"10100011",
		"10100001",
		"10011100",
		"10011011",
		"10011010",
		"10011011",
		"10100001",
		"10100101",
		"10100011",
		"10100000",
		"10100001",
		"10100111",
		"10101101",
		"10110010",
		"10110011",
		"10110001",
		"10101101",
		"01111001",
		"00010110",
		"00001101",
		"00001111",
		"00010001",
		"00010011",
		"00010011",
		"00010100",
		"00010110",
		"00010111",
		"00010111",
		"00011001",
		"00011001",
		"00011001",
		"00011001",
		"00011001",
		"00011010",
		"00011010",
		"00011010",
		"00011011",
		"00011100",
		"00011100",
		"00011111",
		"00011011",
		"00011011",
		"00100011",
		"00101110",
		"00111000",
		"01000101",
		"01011011",
		"01101000",
		"01101100",
		"01011110",
		"01001011",
		"01000111",
		"01000110",
		"01001000",
		"01001000",
		"01001100",
		"01001101",
		"01010011",
		"01010011",
		"01010101",
		"01011101",
		"01011101",
		"01011101",
		"01010111",
		"01000100",
		"00011111",
		"00011100",
		"00010111",
		"00011011",
		"00100000",
		"00100100",
		"00101010",
		"00101101",
		"00101011",
		"00101101",
		"00101000",
		"00100111",
		"00100100",
		"00100001",
		"00100011",
		"00100011",
		"00011011",
		"00010001",
		"00100110",
		"01101110",
		"10111001",
		"11010101",
		"11010101",
		"11010011",
		"11010011",
		"11001000",
		"10101100",
		"10000010",
		"01011000",
		"01100010",
		"01011100",
		"01011011",
		"01101100",
		"01110110",
		"10000111",
		"10011011",
		"10101100",
		"10111111",
		"11001100",
		"11011000",
		"11011011",
		"11011100",
		"11011101",
		"11010111",
		"11010111",
		"11011010",
		"11011010",
		"11010111",
		"11011100",
		"11011010",
		"11010110",
		"11011011",
		"10110001",
		"10010010",
		"10010000",
		"01110101",
		"01011111",
		"01001110",
		"01000100",
		"00111110",
		"01000000",
		"00111110",
		"10001010",
		"11000100",
		"10111110",
		"10111001",
		"10110111",
		"10110010",
		"10110000",
		"10110001",
		"10110001",
		"10110101",
		"10111010",
		"10111101",
		"11000000",
		"10111111",
		"10111111",
		"10111110",
		"10111111",
		"10111110",
		"10111101",
		"10111101",
		"10111110",
		"11000000",
		"10111111",
		"10111110",
		"11000000",
		"10111111",
		"10111110",
		"10111101",
		"10111011",
		"10111100",
		"10111011",
		"10111000",
		"10110011",
		"10110000",
		"10101110",
		"10101110",
		"10101110",
		"10101101",
		"10101001",
		"10010000",
		"01000110",
		"00110011",
		"00111001",
		"00110110",
		"00110010",
		"00101100",
		"00100101",
		"00011111",
		"00011001",
		"00010011",
		"00001110",
		"00001100",
		"00001100",
		"00010000",
		"00010001",
		"00010011",
		"00010101",
		"00010110",
		"00011000",
		"00011010",
		"00011011",
		"00011000",
		"00011100",
		"00100000",
		"00011111",
		"00011010",
		"00011110",
		"00100011",
		"00101111",
		"01000000",
		"01010000",
		"01011100",
		"01001111",
		"00111110",
		"00110111",
		"00111101",
		"01000000",
		"01000011",
		"01001000",
		"01001010",
		"01001101",
		"01010000",
		"01010101",
		"01010100",
		"01010000",
		"01000001",
		"00101111",
		"00011010",
		"00010000",
		"00001110",
		"00010001",
		"00010100",
		"00011001",
		"00100000",
		"00011111",
		"00100011",
		"00100100",
		"00100001",
		"00100010",
		"00011110",
		"00011101",
		"00010111",
		"00010011",
		"00010000",
		"00001111",
		"00001001",
		"00100001",
		"01011111",
		"10111101",
		"11001000",
		"10111001",
		"10111001",
		"10101100",
		"10000101",
		"01110000",
		"01110011",
		"01100101",
		"01011111",
		"01011110",
		"01010111",
		"01101010",
		"01101111",
		"01111101",
		"10001001",
		"10011010",
		"10101101",
		"10111010",
		"11000111",
		"11001011",
		"11001110",
		"11010001",
		"11010011",
		"11010011",
		"11010001",
		"11010110",
		"11011010",
		"11011100",
		"11011100",
		"11011110",
		"11011011",
		"10100100",
		"10000010",
		"10001010",
		"10000011",
		"10001001",
		"01101011",
		"01011111",
		"01010101",
		"01001100",
		"00110101",
		"10001000",
		"10111110",
		"10111000",
		"10110000",
		"10110010",
		"10110110",
		"10111011",
		"10111100",
		"10111100",
		"10111110",
		"10111110",
		"10111101",
		"10111110",
		"10111101",
		"10111110",
		"10111101",
		"10111100",
		"10111100",
		"10111101",
		"10111101",
		"10111100",
		"10111101",
		"10111101",
		"10111100",
		"10111100",
		"10111100",
		"10111101",
		"10111100",
		"10111101",
		"10111110",
		"10111110",
		"10111110",
		"10111101",
		"10111110",
		"10111111",
		"10111101",
		"10111101",
		"10111100",
		"10111010",
		"10110111",
		"10110110",
		"10110110",
		"10110111",
		"10110110",
		"10110101",
		"10110001",
		"10101101",
		"10101000",
		"10100000",
		"10010000",
		"01111100",
		"01100110",
		"01001100",
		"00110100",
		"00011110",
		"00001111",
		"00001011",
		"00001011",
		"00001101",
		"00010001",
		"00010100",
		"00010101",
		"00011000",
		"00011001",
		"00011010",
		"00011101",
		"00011001",
		"00011000",
		"00011101",
		"00100110",
		"00101111",
		"00110100",
		"00110000",
		"00100111",
		"00100101",
		"00101110",
		"00110101",
		"00111001",
		"01000100",
		"01000111",
		"01001100",
		"01001110",
		"01001101",
		"01001001",
		"00111010",
		"00100110",
		"00010100",
		"00001110",
		"00001111",
		"00010000",
		"00010000",
		"00001110",
		"00010001",
		"00011000",
		"00010110",
		"00011011",
		"00011100",
		"00011100",
		"00011100",
		"00011001",
		"00010101",
		"00010110",
		"00010101",
		"00010001",
		"00001110",
		"00001101",
		"00001000",
		"00010111",
		"00110100",
		"00101001",
		"00100011",
		"00111010",
		"01001000",
		"00101010",
		"00010000",
		"00011100",
		"00110000",
		"00111000",
		"00111000",
		"01001011",
		"01101000",
		"01110110",
		"01111111",
		"10000010",
		"10001011",
		"10001101",
		"10100001",
		"10101100",
		"10110011",
		"10110111",
		"10111011",
		"10111110",
		"11000000",
		"10111101",
		"10111011",
		"11000011",
		"11001111",
		"11010100",
		"11010110",
		"11010100",
		"11001011",
		"10010110",
		"01110101",
		"01101111",
		"01100111",
		"01100011",
		"01100110",
		"01100011",
		"01100010",
		"01010001",
		"10000010",
		"10110011",
		"10100110",
		"10100111",
		"10111001",
		"10111101",
		"10111101",
		"10111110",
		"11000000",
		"11000000",
		"11000000",
		"10111111",
		"11000000",
		"10111111",
		"10111111",
		"10111111",
		"10111101",
		"10111100",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111110",
		"10111110",
		"10111110",
		"10111111",
		"10111111",
		"10111111",
		"10111111",
		"10111111",
		"10111110",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111100",
		"10111101",
		"10111110",
		"10111101",
		"10111110",
		"10111100",
		"10111110",
		"10111110",
		"10111111",
		"11000000",
		"11000001",
		"11000010",
		"11000010",
		"11000000",
		"10110111",
		"10101000",
		"10010000",
		"01110010",
		"01011010",
		"01000101",
		"00101111",
		"00011101",
		"00010000",
		"00001110",
		"00010010",
		"00010101",
		"00010111",
		"00010111",
		"00010101",
		"00010010",
		"00010010",
		"00010111",
		"00011110",
		"00011111",
		"00011011",
		"00010111",
		"00011001",
		"00100011",
		"00101101",
		"00111011",
		"01000011",
		"01001010",
		"01000111",
		"00111110",
		"00110001",
		"00011111",
		"00010110",
		"00010010",
		"00010001",
		"00010000",
		"00010000",
		"00010000",
		"00001110",
		"00001101",
		"00001101",
		"00010000",
		"00010001",
		"00010001",
		"00010001",
		"00010001",
		"00010000",
		"00001110",
		"00001111",
		"00001110",
		"00001101",
		"00001100",
		"00001001",
		"00001000",
		"00000110",
		"00000010",
		"00000010",
		"00000010",
		"00000000",
		"00000010",
		"00001111",
		"00011101",
		"00101000",
		"00111010",
		"01000011",
		"01000100",
		"01011001",
		"01011101",
		"01011110",
		"01100001",
		"01100010",
		"01100011",
		"01100000",
		"01100011",
		"01101001",
		"01110010",
		"01110101",
		"01111011",
		"10000011",
		"10000111",
		"10001011",
		"10001101",
		"10010100",
		"10100001",
		"10101001",
		"10101011",
		"10110001",
		"10110010",
		"10010101",
		"10000010",
		"01101100",
		"01011001",
		"01010110",
		"01011000",
		"01011100",
		"01100000",
		"01010110",
		"01110110",
		"10011100",
		"10000010",
		"10100101",
		"10111101",
		"10111101",
		"10111111",
		"11000001",
		"11000001",
		"11000010",
		"11000010",
		"11000010",
		"11000010",
		"11000001",
		"11000001",
		"10111110",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111110",
		"10111101",
		"10111110",
		"10111111",
		"10111110",
		"10111110",
		"10111111",
		"11000000",
		"10111111",
		"10111110",
		"11000000",
		"11000000",
		"10111111",
		"10111111",
		"10111110",
		"10111110",
		"10111111",
		"10111110",
		"10111110",
		"10111111",
		"10111111",
		"10111111",
		"11000000",
		"10111111",
		"10111111",
		"11000000",
		"10111111",
		"11000000",
		"11000000",
		"11000001",
		"11000001",
		"11000000",
		"11000000",
		"10111110",
		"10111111",
		"11000001",
		"11000011",
		"11000000",
		"10111100",
		"10110100",
		"10100100",
		"10000110",
		"01011111",
		"00111000",
		"00011101",
		"00010000",
		"00001110",
		"00010001",
		"00010101",
		"00010110",
		"00010011",
		"00010010",
		"00010011",
		"00010111",
		"00010100",
		"00010100",
		"00011011",
		"00100010",
		"00110011",
		"00111000",
		"00110111",
		"00101111",
		"00100101",
		"00011110",
		"00011000",
		"00010101",
		"00010100",
		"00010101",
		"00010100",
		"00010000",
		"00010000",
		"00010000",
		"00010000",
		"00001111",
		"00001111",
		"00001101",
		"00001101",
		"00001110",
		"00001101",
		"00001100",
		"00001101",
		"00001100",
		"00001100",
		"00001010",
		"00001001",
		"00001001",
		"00000111",
		"00000101",
		"00000110",
		"00001110",
		"00011010",
		"00110010",
		"01001110",
		"01011100",
		"01011111",
		"01100000",
		"01011101",
		"01011011",
		"01011100",
		"01011001",
		"01011000",
		"01011000",
		"01011001",
		"01011011",
		"01011100",
		"01011010",
		"01011000",
		"01010111",
		"01010101",
		"01010100",
		"01010001",
		"01001101",
		"01001100",
		"01001101",
		"01001101",
		"01001101",
		"01010001",
		"01010100",
		"01010110",
		"01011000",
		"01011010",
		"01011111",
		"01100010",
		"01100000",
		"01011011",
		"01100000",
		"01100011",
		"01011011",
		"01010101",
		"01001010",
		"01010000",
		"01010111",
		"01010001",
		"10101100",
		"11000001",
		"11000000",
		"11000011",
		"11000100",
		"11000100",
		"11000101",
		"11000110",
		"11000110",
		"11000101",
		"11000100",
		"11000011",
		"11000001",
		"11000001",
		"11000000",
		"11000000",
		"10111111",
		"10111111",
		"11000000",
		"11000000",
		"10111111",
		"11000001",
		"11000010",
		"11000001",
		"11000001",
		"11000001",
		"11000000",
		"11000000",
		"11000001",
		"11000000",
		"11000001",
		"11000000",
		"10111111",
		"11000000",
		"11000001",
		"11000010",
		"11000010",
		"11000010",
		"11000001",
		"11000000",
		"11000000",
		"11000000",
		"11000011",
		"11000101",
		"11000110",
		"11001000",
		"11000111",
		"11000101",
		"11000101",
		"11000100",
		"11000011",
		"11000011",
		"11000011",
		"11000011",
		"11000010",
		"11000011",
		"11000010",
		"11000010",
		"11000100",
		"11000100",
		"10111011",
		"10100101",
		"10000101",
		"01011111",
		"00110110",
		"00011010",
		"00011100",
		"00011011",
		"00011011",
		"00011010",
		"00011001",
		"00011100",
		"00100100",
		"00100111",
		"00101110",
		"00110100",
		"00110110",
		"00110111",
		"00110110",
		"00110110",
		"00110111",
		"00111001",
		"00111100",
		"00111101",
		"00111111",
		"00111011",
		"00110101",
		"00101110",
		"00101010",
		"00100101",
		"00100001",
		"00011100",
		"00010111",
		"00010110",
		"00010100",
		"00010001",
		"00001110",
		"00001101",
		"00001100",
		"00001011",
		"00001010",
		"00000111",
		"00000111",
		"00001101",
		"00011101",
		"00110001",
		"01000101",
		"01001110",
		"01010111",
		"01011001",
		"01010111",
		"01010111",
		"01010101",
		"01010011",
		"01010100",
		"01010100",
		"01010000",
		"01010010",
		"01010010",
		"01010011",
		"01010100",
		"01010011",
		"01010001",
		"01010100",
		"01010110",
		"01010100",
		"01010101",
		"01010111",
		"01011000",
		"01010110",
		"01011000",
		"01011011",
		"01011011",
		"01011000",
		"01011010",
		"01011010",
		"01011001",
		"01011010",
		"01011101",
		"01011111",
		"01100110",
		"01111011",
		"10011011",
		"10100100",
		"10010000",
		"10000011",
		"01110111",
		"00101111",
		"00111100",
		"10000101",
		"10101100",
		"10111100",
		"11000001",
		"11000011",
		"11000100",
		"11000100",
		"11000101",
		"11000110",
		"11000111",
		"11001000",
		"11000101",
		"11000101",
		"11000011",
		"11000010",
		"11000010",
		"11000000",
		"11000000",
		"11000001",
		"11000001",
		"11000000",
		"10111111",
		"11000001",
		"11000001",
		"11000010",
		"11000011",
		"11001000",
		"11000010",
		"11000000",
		"11000001",
		"11000001",
		"11000000",
		"11000001",
		"11000001",
		"11000010",
		"11000111",
		"11001001",
		"11000111",
		"11001000",
		"11000111",
		"11000100",
		"11000110",
		"11001001",
		"11001100",
		"11001111",
		"11010001",
		"11010011",
		"11010001",
		"11010001",
		"11010001",
		"11010010",
		"11010010",
		"11010000",
		"11001110",
		"11001111",
		"11001101",
		"11001100",
		"11001010",
		"11000111",
		"11000110",
		"11000110",
		"11000101",
		"11000111",
		"11001010",
		"11001011",
		"10111110",
		"01110011",
		"00101001",
		"00110000",
		"00110111",
		"00111111",
		"01000000",
		"01000110",
		"01001000",
		"01000010",
		"01000000",
		"01000110",
		"01001100",
		"01001111",
		"01010000",
		"01010001",
		"01010100",
		"01010111",
		"01011100",
		"01011101",
		"01100000",
		"01011110",
		"01100000",
		"01011111",
		"01100000",
		"01011101",
		"01011010",
		"01010111",
		"01010101",
		"01010011",
		"01001111",
		"01000111",
		"00111110",
		"00111001",
		"00111010",
		"00111010",
		"00111011",
		"01000011",
		"01010010",
		"01011110",
		"01100110",
		"01011101",
		"01001111",
		"01001101",
		"01010010",
		"01010111",
		"01011000",
		"01011000",
		"01010111",
		"01010101",
		"01010001",
		"01010001",
		"01001111",
		"01001110",
		"01001101",
		"01010001",
		"01010011",
		"01000001",
		"01000110",
		"01001010",
		"01001010",
		"01001011",
		"01001110",
		"01001111",
		"01001111",
		"01010000",
		"01010100",
		"01010101",
		"01010110",
		"01010110",
		"01010111",
		"01011010",
		"01011101",
		"01100001",
		"01100111",
		"01101010",
		"01110110",
		"10011001",
		"10111000",
		"10110111",
		"10111111",
		"10101101",
		"10100110",
		"00111001",
		"01101111",
		"10101000",
		"10010010",
		"10101010",
		"10111110",
		"11000000",
		"11000010",
		"11000010",
		"11000011",
		"11000100",
		"11000101",
		"11000100",
		"11000010",
		"11000010",
		"11000010",
		"11000010",
		"11000001",
		"10111111",
		"10111111",
		"11000001",
		"11000000",
		"11000000",
		"11000000",
		"11000001",
		"11000000",
		"11000010",
		"11000101",
		"11001010",
		"11000110",
		"10111110",
		"10111111",
		"11000001",
		"11000001",
		"11000110",
		"11001010",
		"11001001",
		"11001010",
		"11001101",
		"11001011",
		"11001111",
		"11010010",
		"11010101",
		"11010101",
		"11010011",
		"11001111",
		"11001010",
		"11000101",
		"11000000",
		"11000000",
		"10111111",
		"11000001",
		"11000110",
		"11001001",
		"11001001",
		"11001001",
		"11001010",
		"11001100",
		"11010001",
		"11010010",
		"11010010",
		"11001111",
		"11001100",
		"11001111",
		"11010000",
		"11010000",
		"11001101",
		"11001000",
		"10100100",
		"01001100",
		"01000111",
		"01000010",
		"00111101",
		"00110010",
		"00110001",
		"00110110",
		"00111101",
		"01000100",
		"01001001",
		"01001101",
		"01001111",
		"01010001",
		"01010100",
		"01010111",
		"01010100",
		"01010100",
		"01010110",
		"01011000",
		"01011001",
		"01011010",
		"01011011",
		"01011011",
		"01011001",
		"01011000",
		"01011001",
		"01011001",
		"01011000",
		"01010110",
		"01010110",
		"01010110",
		"01010101",
		"01010110",
		"01011001",
		"01100001",
		"01110000",
		"10000100",
		"10001011",
		"10011001",
		"10101001",
		"10011100",
		"01111101",
		"01011001",
		"01001110",
		"01010111",
		"01011010",
		"01011000",
		"01010110",
		"01010110",
		"01010011",
		"01010010",
		"01001111",
		"01010010",
		"01010110",
		"01010011",
		"01001011",
		"01111100",
		"01011001",
		"01001101",
		"01001111",
		"01010000",
		"01010010",
		"01010011",
		"01010101",
		"01011000",
		"01011010",
		"01011010",
		"01010111",
		"01011010",
		"01011100",
		"01011110",
		"01100100",
		"01101101",
		"10001010",
		"10010100",
		"10111101",
		"11000101",
		"10000110",
		"10110010",
		"10111011",
		"10110000",
		"01100110",
		"10000101",
		"10100000",
		"10001100",
		"10100011",
		"10111110",
		"10111111",
		"11000001",
		"11000001",
		"11000001",
		"11000010",
		"11000011",
		"11000011",
		"11000000",
		"11000000",
		"11000000",
		"11000000",
		"10111110",
		"10111101",
		"10111101",
		"10111101",
		"10111101",
		"10111110",
		"10111111",
		"11000000",
		"11000010",
		"11000100",
		"11000101",
		"11001010",
		"11001001",
		"11000000",
		"11000000",
		"11000011",
		"11000011",
		"11001010",
		"11010001",
		"11001100",
		"11000101",
		"11000111",
		"11001010",
		"11001000",
		"11000000",
		"10111000",
		"10110011",
		"10101101",
		"10101100",
		"10101011",
		"10101101",
		"10110000",
		"10110100",
		"10110110",
		"10111011",
		"10111110",
		"10111111",
		"11000000",
		"11000000",
		"10111111",
		"10111111",
		"11000000",
		"10111101",
		"10111100",
		"10111011",
		"10111010",
		"10111000",
		"10111000",
		"10110110",
		"10110101",
		"10110101",
		"10110011",
		"10101111",
		"10101111",
		"10101011",
		"10100001",
		"10001011",
		"01101001",
		"01001100",
		"01000010",
		"00111110",
		"00111100",
		"01000100",
		"01010000",
		"01011000",
		"01011100",
		"01011111",
		"01011100",
		"01011001",
		"01011001",
		"01011001",
		"01011010",
		"01011100",
		"01011100",
		"01011000",
		"01011001",
		"01011001",
		"01010101",
		"01010100",
		"01010001",
		"01010000",
		"01010001",
		"01010010",
		"01011000",
		"01011101",
		"01100100",
		"01101011",
		"01111010",
		"10001011",
		"10011010",
		"10011110",
		"10101001",
		"11000001",
		"10101001",
		"10010101",
		"01011100",
		"01000110",
		"01001011",
		"01001110",
		"01010000",
		"01010010",
		"01010010",
		"01010011",
		"01010101",
		"01010111",
		"01010101",
		"01001011",
		"01011100",
		"10010011",
		"10010000",
		"01010101",
		"01010101",
		"01010111",
		"01010111",
		"01011000",
		"01011000",
		"01011011",
		"01011101",
		"01011100",
		"01011100",
		"01011111",
		"01011110",
		"01100100",
		"01101101",
		"01110111",
		"10010110",
		"10101101",
		"10111111",
		"10111110",
		"10110101",
		"10111000",
		"11000000",
		"11000111",
		"01011011",
		"01110001",
		"10001101",
		"10101000",
		"10101111",
		"10111101",
		"10111110",
		"11000000",
		"10111111",
		"10111111",
		"10111111",
		"11000010",
		"11000011",
		"11000001",
		"11000001",
		"11000010",
		"11000001",
		"11000000",
		"11000000",
		"11000000",
		"10111110",
		"10111110",
		"10111110",
		"11000000",
		"11000100",
		"11000100",
		"11000100",
		"11000100",
		"11000110",
		"11000110",
		"11000001",
		"11000000",
		"11000000",
		"10111110",
		"10111100",
		"10111101",
		"10111101",
		"10111010",
		"10111001",
		"10110000",
		"10101000",
		"10100110",
		"10101010",
		"10101110",
		"10110010",
		"10110101",
		"10110111",
		"10111001",
		"10111010",
		"10111010",
		"10111101",
		"11000010",
		"11000011",
		"11000100",
		"11000101",
		"11000110",
		"11001000",
		"11001010",
		"11001001",
		"11000111",
		"11000101",
		"11000011",
		"11000001",
		"11000010",
		"11000011",
		"11000101",
		"11000110",
		"11000101",
		"11000101",
		"11000111",
		"11000110",
		"11000111",
		"11001010",
		"11001100",
		"11001101",
		"11001001",
		"10111011",
		"10101001",
		"10001101",
		"01100001",
		"01000101",
		"01001001",
		"01010000",
		"01011000",
		"01011111",
		"01100011",
		"01100100",
		"01100100",
		"01100000",
		"01011111",
		"01100000",
		"01011101",
		"01011101",
		"01011100",
		"01011000",
		"01010110",
		"01010110",
		"01011000",
		"01011001",
		"01011110",
		"01100111",
		"01110001",
		"01110100",
		"10000000",
		"10010011",
		"10101010",
		"11000010",
		"10100110",
		"10010001",
		"10100101",
		"10101001",
		"10101001",
		"10001001",
		"01001111",
		"01000111",
		"01001011",
		"01001101",
		"01001111",
		"01001111",
		"01010001",
		"01010001",
		"01001010",
		"00110110",
		"01011001",
		"10011011",
		"10001111",
		"01100001",
		"01010100",
		"01010101",
		"01010101",
		"01010010",
		"01010000",
		"01010011",
		"01010111",
		"01011000",
		"01011100",
		"01011101",
		"01011101",
		"01100010",
		"01101101",
		"01101111",
		"10000011",
		"10011001",
		"10111101",
		"11010000",
		"10101110",
		"11000011",
		"11001010",
		"11000111",
		"11000000"
			);

begin

addr_1 <= addr;
addr_2 <= addr + 1;
addr_3 <= addr + 299;
addr_4 <= addr + 300;

process(clk)
begin
  if(rising_edge(clk)) then
    if (rst = '1') then
      data_o_1 <= "00000000";
    else
      data_o_1 <= rom(addr);
      data_o_2 <= rom(addr_2);
      data_o_3 <= rom(addr_3);
      data_o_4 <= rom(addr_4);
    end if;
  end if;
end process;
end arch;
