--Engineer     : Navdeep Dahiya
--Date         : 11/15/2018
--Name of file : block_rom.vhd
--Description  : module ROM as block rom

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity blk_rom is
  port (
	-- input side
	clk	: in std_logic;
	rst	: in std_logic;
	addr	: in integer range 0 to 255; -- address bits
	--output side
	data_o	: out std_logic_vector(7 downto 0)
	);
end blk_rom;

architecture arch of blk_rom is

type rom_t is array(0 to 255) of std_logic_vector(7 downto 0);

signal rom : rom_t := (
		"00011110",
		"00111010",
		"00111110",
		"01000000",
		"01000001",
		"00111001",
		"00110111",
		"00111000",
		"00111001",
		"00111000",
		"01001010",
		"01001000",
		"01001001",
		"01001100",
		"01001001",
		"01001111",
		"00100101",
		"01110111",
		"01110010",
		"01110011",
		"01110011",
		"01110100",
		"01101111",
		"01101010",
		"01110001",
		"01101011",
		"01101101",
		"01101100",
		"01110000",
		"01101111",
		"01101100",
		"01101000",
		"00100110",
		"01111001",
		"01110011",
		"01101101",
		"01110000",
		"01101110",
		"01110010",
		"01101000",
		"01110001",
		"01110010",
		"01101111",
		"01101111",
		"01101110",
		"01110001",
		"01100011",
		"01101110",
		"00100101",
		"01101100",
		"01111001",
		"01101101",
		"01110010",
		"01110001",
		"01101001",
		"01101101",
		"01100111",
		"01101010",
		"01101101",
		"01101001",
		"01110110",
		"01110000",
		"01100010",
		"01101110",
		"00100110",
		"01110011",
		"01111100",
		"01110110",
		"01101110",
		"01110110",
		"01101010",
		"01110000",
		"01101010",
		"01101111",
		"01110000",
		"01101110",
		"01110010",
		"01101001",
		"01101010",
		"01100110",
		"00100101",
		"01110010",
		"01110110",
		"01101010",
		"01110001",
		"01101101",
		"01110001",
		"01101111",
		"01101100",
		"01101101",
		"01100101",
		"01101011",
		"01110010",
		"01110001",
		"01101100",
		"01101000",
		"00100100",
		"01101110",
		"01101011",
		"01110001",
		"01100111",
		"01110010",
		"01101110",
		"01110000",
		"01101010",
		"01101000",
		"01101101",
		"01110010",
		"01110010",
		"01101100",
		"01110001",
		"01101000",
		"00100100",
		"01101110",
		"01110011",
		"01100111",
		"01101110",
		"01110001",
		"01110001",
		"01100110",
		"01110000",
		"01101101",
		"01101010",
		"01110001",
		"01110010",
		"01110000",
		"01101101",
		"01110001",
		"00100011",
		"01100010",
		"01101101",
		"01110100",
		"01101011",
		"01110001",
		"01101011",
		"01101110",
		"01101001",
		"01101011",
		"01110001",
		"01100110",
		"01110000",
		"01101101",
		"01110001",
		"01110011",
		"00100000",
		"01101101",
		"01110100",
		"01101001",
		"01101111",
		"01110001",
		"01110101",
		"01101011",
		"01100110",
		"01110001",
		"01101100",
		"01101101",
		"01101011",
		"01110110",
		"01101110",
		"01101110",
		"00011000",
		"01110000",
		"01101100",
		"01110011",
		"01100110",
		"01101101",
		"01110000",
		"01100101",
		"01100111",
		"01101001",
		"01101010",
		"01101000",
		"01101000",
		"01101100",
		"01101101",
		"01101011",
		"00010110",
		"01100111",
		"01110001",
		"01101111",
		"01101100",
		"01110010",
		"01101110",
		"01101011",
		"01101011",
		"01101010",
		"01101001",
		"01110000",
		"01100110",
		"01110001",
		"01100100",
		"01101011",
		"00010011",
		"01101001",
		"01101100",
		"01101110",
		"01100100",
		"01101101",
		"01011101",
		"01100011",
		"01100011",
		"01101101",
		"01101111",
		"01101001",
		"01101110",
		"01100100",
		"01110000",
		"01100101",
		"00010010",
		"01100101",
		"01101100",
		"01110000",
		"01100001",
		"01101011",
		"01100111",
		"01101010",
		"01011011",
		"01101001",
		"01101011",
		"01100111",
		"01100101",
		"01100111",
		"01101010",
		"01100011",
		"00010101",
		"01110000",
		"01101100",
		"01101001",
		"01101010",
		"01100100",
		"01100010",
		"01100000",
		"01100011",
		"01101100",
		"01100100",
		"01101001",
		"01100101",
		"01101111",
		"01100101",
		"01100101",
		"00010011",
		"01101000",
		"01101100",
		"01101011",
		"01100000",
		"01101011",
		"01101001",
		"01101000",
		"01100111",
		"01110001",
		"01101110",
		"01101011",
		"01101101",
		"01101111",
		"01110101",
		"01101011"
			);

begin

process(clk)
begin
  if(rising_edge(clk)) then
    if (rst = '1') then
      data_o <= "00000000";
    else
      data_o <= rom(addr);
    end if;
  end if;
end process;
end arch;
